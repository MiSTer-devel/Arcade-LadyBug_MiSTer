library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"B8",X"CA",X"03",X"21",X"11",X"05",X"00",X"DD",X"19",X"C3",X"F5",X"1F",X"21",X"5F",X"60",X"CB",
		X"4E",X"28",X"20",X"21",X"02",X"90",X"CB",X"6E",X"28",X"19",X"4F",X"3A",X"65",X"60",X"FE",X"00",
		X"79",X"28",X"10",X"DD",X"4E",X"02",X"3E",X"FE",X"91",X"4F",X"DD",X"56",X"01",X"3E",X"AE",X"92",
		X"C3",X"39",X"20",X"DD",X"7E",X"01",X"DD",X"4E",X"02",X"DD",X"56",X"00",X"CB",X"3A",X"CB",X"3A",
		X"CB",X"3A",X"CB",X"3A",X"CD",X"A8",X"1F",X"D5",X"16",X"00",X"FD",X"21",X"4E",X"60",X"FD",X"19",
		X"F5",X"FD",X"7E",X"00",X"FD",X"34",X"00",X"C5",X"43",X"04",X"FD",X"21",X"80",X"70",X"11",X"40",
		X"00",X"FD",X"19",X"10",X"FC",X"CB",X"27",X"CB",X"27",X"5F",X"FD",X"19",X"C1",X"79",X"D6",X"07",
		X"FD",X"77",X"03",X"F1",X"E6",X"0F",X"D1",X"1E",X"00",X"CB",X"52",X"20",X"06",X"CB",X"42",X"28",
		X"06",X"CB",X"E7",X"1C",X"C3",X"8D",X"20",X"CB",X"5A",X"20",X"02",X"CB",X"EF",X"21",X"5F",X"60",
		X"CB",X"4E",X"28",X"2A",X"21",X"02",X"90",X"CB",X"6E",X"28",X"23",X"32",X"C8",X"61",X"3A",X"65",
		X"60",X"FE",X"00",X"3A",X"C8",X"61",X"28",X"16",X"CB",X"67",X"20",X"05",X"CB",X"E7",X"C3",X"B3",
		X"20",X"CB",X"A7",X"CB",X"6F",X"20",X"05",X"CB",X"EF",X"C3",X"BE",X"20",X"CB",X"AF",X"F6",X"C0",
		X"FD",X"77",X"00",X"DD",X"7E",X"03",X"DD",X"CB",X"04",X"66",X"20",X"2B",X"FE",X"D8",X"30",X"27",
		X"08",X"AF",X"BB",X"20",X"06",X"08",X"C6",X"0C",X"C3",X"DC",X"20",X"08",X"08",X"3A",X"5A",X"60",
		X"E6",X"03",X"CB",X"47",X"28",X"05",X"16",X"04",X"C3",X"F1",X"20",X"FE",X"02",X"20",X"07",X"16",
		X"08",X"08",X"82",X"C3",X"F7",X"20",X"08",X"FD",X"77",X"01",X"DD",X"7E",X"04",X"FD",X"77",X"02",
		X"C3",X"FD",X"1F",X"21",X"C0",X"70",X"06",X"0B",X"DD",X"21",X"4E",X"60",X"DD",X"7E",X"00",X"E5",
		X"CB",X"27",X"CB",X"27",X"5F",X"16",X"00",X"19",X"72",X"E5",X"D1",X"7B",X"D1",X"D5",X"93",X"FE",
		X"20",X"30",X"0D",X"FD",X"E1",X"FD",X"E5",X"11",X"20",X"00",X"FD",X"19",X"AF",X"FD",X"77",X"00",
		X"11",X"40",X"00",X"DD",X"23",X"E1",X"19",X"10",X"D3",X"21",X"01",X"90",X"CB",X"7E",X"C2",X"3C",
		X"21",X"DD",X"E1",X"C9",X"3E",X"00",X"06",X"16",X"21",X"A6",X"D4",X"11",X"20",X"00",X"C5",X"06",
		X"16",X"E5",X"77",X"23",X"10",X"FC",X"E1",X"C1",X"19",X"10",X"F3",X"C9",X"DD",X"21",X"E7",X"D0",
		X"3E",X"32",X"11",X"20",X"00",X"DD",X"77",X"01",X"DD",X"77",X"05",X"DD",X"77",X"07",X"DD",X"77",
		X"08",X"DD",X"77",X"11",X"3D",X"DD",X"77",X"04",X"DD",X"77",X"0A",X"DD",X"77",X"0C",X"3D",X"DD",
		X"77",X"02",X"3C",X"DD",X"19",X"DD",X"77",X"02",X"DD",X"77",X"04",X"DD",X"77",X"0A",X"DD",X"77",
		X"0C",X"DD",X"77",X"10",X"DD",X"19",X"3C",X"DD",X"77",X"09",X"DD",X"77",X"0A",X"DD",X"77",X"0D",
		X"3C",X"DD",X"77",X"04",X"DD",X"77",X"0C",X"DD",X"77",X"10",X"DD",X"19",X"3D",X"3D",X"DD",X"77",
		X"02",X"DD",X"19",X"DD",X"77",X"00",X"3C",X"DD",X"77",X"05",X"DD",X"77",X"0B",X"DD",X"77",X"11",
		X"DD",X"77",X"12",X"3C",X"DD",X"77",X"04",X"DD",X"19",X"3D",X"3D",X"DD",X"77",X"00",X"DD",X"19",
		X"3C",X"DD",X"77",X"09",X"DD",X"77",X"0A",X"3C",X"DD",X"77",X"00",X"DD",X"19",X"3D",X"3D",X"DD",
		X"77",X"04",X"DD",X"77",X"0E",X"DD",X"77",X"12",X"DD",X"19",X"DD",X"77",X"08",X"3C",X"DD",X"77",
		X"01",X"DD",X"77",X"02",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"09",X"DD",X"77",X"0A",
		X"DD",X"77",X"0D",X"DD",X"77",X"0E",X"DD",X"77",X"11",X"DD",X"77",X"12",X"3C",X"DD",X"77",X"00",
		X"DD",X"77",X"04",X"DD",X"77",X"0C",X"DD",X"77",X"10",X"DD",X"19",X"3D",X"3D",X"DD",X"77",X"08",
		X"DD",X"19",X"3D",X"DD",X"77",X"0E",X"DD",X"77",X"12",X"3C",X"DD",X"77",X"04",X"3C",X"DD",X"77",
		X"01",X"DD",X"77",X"05",X"DD",X"77",X"09",X"DD",X"77",X"0A",X"DD",X"77",X"0D",X"DD",X"77",X"11",
		X"3C",X"DD",X"77",X"00",X"DD",X"77",X"08",X"DD",X"19",X"3D",X"3D",X"DD",X"77",X"04",X"DD",X"77",
		X"0E",X"DD",X"77",X"12",X"DD",X"19",X"DD",X"77",X"00",X"3C",X"DD",X"77",X"09",X"DD",X"77",X"0A",
		X"DD",X"19",X"3D",X"DD",X"77",X"00",X"DD",X"19",X"DD",X"77",X"02",X"3C",X"DD",X"77",X"05",X"DD",
		X"77",X"0B",X"DD",X"77",X"0C",X"DD",X"77",X"11",X"3C",X"DD",X"77",X"04",X"DD",X"19",X"3D",X"3D",
		X"DD",X"77",X"02",X"DD",X"19",X"DD",X"77",X"04",X"DD",X"77",X"0C",X"DD",X"77",X"10",X"3C",X"DD",
		X"77",X"09",X"DD",X"77",X"0D",X"3D",X"3D",X"DD",X"77",X"0A",X"DD",X"19",X"3C",X"DD",X"77",X"02",
		X"DD",X"77",X"04",X"DD",X"77",X"0A",X"DD",X"77",X"0C",X"DD",X"77",X"10",X"DD",X"19",X"3C",X"DD",
		X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"77",
		X"08",X"DD",X"77",X"11",X"DD",X"77",X"12",X"3C",X"DD",X"77",X"00",X"DD",X"77",X"04",X"DD",X"77",
		X"0A",X"DD",X"77",X"0C",X"C9",X"E5",X"C5",X"06",X"FF",X"C5",X"06",X"FF",X"C5",X"06",X"FF",X"00",
		X"10",X"FD",X"C1",X"10",X"F7",X"C1",X"10",X"F1",X"C1",X"E1",X"C9",X"E5",X"C5",X"E5",X"FE",X"04",
		X"38",X"10",X"CB",X"47",X"28",X"06",X"FD",X"21",X"F0",X"0C",X"18",X"52",X"FD",X"21",X"E7",X"0C",
		X"18",X"4C",X"0E",X"00",X"CB",X"47",X"28",X"24",X"11",X"E1",X"FF",X"19",X"08",X"7E",X"FE",X"E5",
		X"20",X"02",X"CB",X"C1",X"11",X"3E",X"00",X"19",X"7E",X"FE",X"E5",X"20",X"02",X"CB",X"D9",X"F5",
		X"79",X"32",X"8E",X"60",X"F1",X"08",X"FD",X"21",X"DE",X"0C",X"18",X"22",X"11",X"21",X"00",X"19",
		X"08",X"7E",X"FE",X"E5",X"20",X"02",X"CB",X"C9",X"11",X"BE",X"FF",X"19",X"7E",X"FE",X"E5",X"20",
		X"02",X"CB",X"D1",X"F5",X"79",X"32",X"8E",X"60",X"F1",X"08",X"FD",X"21",X"D5",X"0C",X"CD",X"0F",
		X"24",X"E1",X"0E",X"00",X"08",X"CB",X"3A",X"CB",X"1B",X"D2",X"DF",X"23",X"79",X"FE",X"00",X"20",
		X"05",X"CD",X"D9",X"24",X"18",X"79",X"FE",X"04",X"20",X"05",X"CD",X"8B",X"24",X"18",X"70",X"CD",
		X"23",X"24",X"D5",X"FD",X"E5",X"16",X"00",X"3D",X"FE",X"04",X"38",X"01",X"3D",X"5F",X"FD",X"19",
		X"FD",X"7E",X"00",X"FD",X"E1",X"D1",X"FE",X"01",X"20",X"40",X"E5",X"21",X"8E",X"60",X"79",X"FE",
		X"03",X"20",X"06",X"CB",X"4E",X"28",X"18",X"18",X"1A",X"30",X"06",X"CB",X"46",X"28",X"10",X"18",
		X"12",X"FE",X"08",X"20",X"06",X"CB",X"56",X"28",X"06",X"18",X"08",X"CB",X"5E",X"20",X"04",X"3E",
		X"FF",X"18",X"14",X"3E",X"E5",X"F5",X"3E",X"02",X"DD",X"E5",X"D5",X"11",X"00",X"04",X"DD",X"19",
		X"DD",X"77",X"00",X"D1",X"DD",X"E1",X"F1",X"E1",X"18",X"12",X"F5",X"3E",X"00",X"DD",X"E5",X"D5",
		X"11",X"00",X"04",X"DD",X"19",X"DD",X"77",X"00",X"D1",X"DD",X"E1",X"F1",X"DD",X"77",X"00",X"79",
		X"FE",X"0A",X"28",X"05",X"0C",X"08",X"C3",X"54",X"23",X"08",X"FE",X"04",X"38",X"0D",X"3E",X"00",
		X"32",X"8E",X"60",X"32",X"90",X"60",X"32",X"8F",X"60",X"18",X"11",X"3E",X"09",X"32",X"8F",X"60",
		X"3E",X"01",X"32",X"90",X"60",X"E5",X"21",X"00",X"60",X"CB",X"C6",X"E1",X"C1",X"E1",X"C9",X"F5",
		X"CB",X"27",X"5F",X"16",X"00",X"DD",X"21",X"F9",X"0C",X"DD",X"19",X"DD",X"56",X"00",X"DD",X"5E",
		X"01",X"F1",X"C9",X"D5",X"E5",X"DD",X"E1",X"FE",X"06",X"28",X"3C",X"FE",X"02",X"20",X"04",X"DD",
		X"23",X"18",X"34",X"30",X"07",X"11",X"E1",X"FF",X"DD",X"19",X"18",X"2B",X"FE",X"05",X"20",X"05",
		X"11",X"E0",X"FF",X"18",X"F3",X"30",X"05",X"11",X"21",X"00",X"18",X"EC",X"FE",X"08",X"20",X"05",
		X"11",X"DF",X"FF",X"18",X"E3",X"30",X"05",X"11",X"20",X"00",X"18",X"DC",X"FE",X"09",X"28",X"05",
		X"11",X"1F",X"00",X"18",X"D3",X"DD",X"2B",X"D1",X"C9",X"DD",X"21",X"09",X"0D",X"78",X"3D",X"16",
		X"00",X"5F",X"DD",X"19",X"DD",X"56",X"00",X"79",X"FE",X"00",X"28",X"0B",X"CB",X"3A",X"CB",X"3A",
		X"CB",X"3A",X"CB",X"3A",X"7A",X"18",X"03",X"7A",X"E6",X"0F",X"C9",X"D5",X"E5",X"11",X"C0",X"FF",
		X"19",X"CD",X"69",X"24",X"FE",X"02",X"20",X"0D",X"08",X"FE",X"04",X"38",X"04",X"36",X"34",X"18",
		X"34",X"36",X"33",X"18",X"30",X"30",X"0D",X"08",X"FE",X"04",X"38",X"04",X"36",X"38",X"18",X"25",
		X"36",X"32",X"18",X"21",X"08",X"FE",X"04",X"38",X"0E",X"08",X"7E",X"FE",X"3B",X"20",X"04",X"36",
		X"3A",X"18",X"13",X"36",X"34",X"18",X"0F",X"08",X"7E",X"FE",X"3A",X"20",X"04",X"36",X"3B",X"18",
		X"05",X"36",X"33",X"18",X"01",X"08",X"E1",X"D1",X"C9",X"D5",X"E5",X"23",X"23",X"CD",X"69",X"24",
		X"FE",X"02",X"20",X"0D",X"08",X"FE",X"04",X"38",X"04",X"36",X"3B",X"18",X"34",X"36",X"33",X"18",
		X"30",X"30",X"0D",X"08",X"FE",X"04",X"38",X"04",X"36",X"3C",X"18",X"25",X"36",X"31",X"18",X"21",
		X"08",X"FE",X"04",X"38",X"0E",X"08",X"7E",X"FE",X"34",X"20",X"04",X"36",X"3A",X"18",X"13",X"36",
		X"3B",X"18",X"0F",X"08",X"7E",X"FE",X"3A",X"20",X"04",X"36",X"34",X"18",X"05",X"36",X"33",X"18",
		X"01",X"08",X"E1",X"D1",X"C9",X"CD",X"06",X"2B",X"CD",X"BA",X"1A",X"CD",X"55",X"17",X"CD",X"3E",
		X"25",X"CD",X"07",X"26",X"CD",X"1D",X"27",X"CD",X"CB",X"27",X"CD",X"26",X"28",X"C9",X"06",X"10",
		X"21",X"1E",X"D1",X"DD",X"21",X"D7",X"2E",X"0E",X"06",X"CD",X"B3",X"27",X"21",X"DC",X"D0",X"06",
		X"01",X"E5",X"78",X"FE",X"01",X"28",X"08",X"0E",X"03",X"CD",X"B1",X"25",X"77",X"18",X"07",X"0E",
		X"07",X"CD",X"B1",X"25",X"36",X"1D",X"11",X"20",X"00",X"19",X"DD",X"21",X"CF",X"2E",X"FE",X"05",
		X"30",X"08",X"3D",X"CB",X"27",X"16",X"00",X"5F",X"18",X"03",X"11",X"06",X"00",X"DD",X"19",X"CD",
		X"B1",X"25",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"D5",X"11",X"20",X"00",X"19",X"D1",X"CD",X"B1",
		X"25",X"DD",X"7E",X"00",X"77",X"D5",X"11",X"40",X"00",X"19",X"D1",X"CD",X"BD",X"25",X"E1",X"04",
		X"78",X"FE",X"0A",X"30",X"0B",X"FE",X"02",X"20",X"04",X"2B",X"2B",X"18",X"A4",X"2B",X"18",X"A1",
		X"C9",X"F5",X"E5",X"D5",X"11",X"00",X"04",X"19",X"71",X"D1",X"E1",X"F1",X"C9",X"78",X"DD",X"21",
		X"80",X"D3",X"3D",X"CB",X"27",X"CB",X"27",X"57",X"CB",X"27",X"82",X"5F",X"16",X"00",X"DD",X"19",
		X"C5",X"06",X"0C",X"11",X"00",X"04",X"E5",X"19",X"71",X"E1",X"DD",X"7E",X"00",X"77",X"D5",X"11",
		X"20",X"00",X"19",X"DD",X"23",X"D1",X"10",X"EE",X"06",X"06",X"79",X"E5",X"19",X"CD",X"7D",X"1E",
		X"E1",X"C1",X"DD",X"21",X"73",X"60",X"78",X"C5",X"3D",X"47",X"CB",X"27",X"80",X"C1",X"5F",X"16",
		X"00",X"DD",X"19",X"CD",X"06",X"1E",X"C9",X"21",X"AC",X"D4",X"3E",X"02",X"0E",X"07",X"11",X"20",
		X"00",X"E5",X"06",X"17",X"77",X"19",X"10",X"FC",X"E1",X"23",X"0D",X"20",X"F4",X"21",X"50",X"D7",
		X"3E",X"07",X"77",X"23",X"77",X"19",X"77",X"2B",X"77",X"21",X"B1",X"D0",X"3E",X"AA",X"CD",X"F6",
		X"26",X"2B",X"2B",X"36",X"BC",X"2B",X"3E",X"B4",X"77",X"3C",X"19",X"77",X"19",X"77",X"19",X"E5",
		X"36",X"A5",X"19",X"36",X"A6",X"E1",X"23",X"3E",X"A7",X"CD",X"07",X"27",X"2B",X"A7",X"ED",X"52",
		X"3E",X"A4",X"CD",X"07",X"27",X"21",X"6F",X"D1",X"36",X"A7",X"19",X"36",X"A8",X"21",X"B1",X"D1",
		X"3E",X"AA",X"CD",X"F6",X"26",X"2B",X"2B",X"E5",X"3E",X"B1",X"CD",X"07",X"27",X"E1",X"2B",X"3E",
		X"A4",X"CD",X"07",X"27",X"21",X"0F",X"D2",X"36",X"BD",X"2B",X"36",X"BF",X"2B",X"36",X"AD",X"A7",
		X"ED",X"52",X"36",X"AE",X"2B",X"3E",X"BB",X"CD",X"11",X"27",X"21",X"51",X"D2",X"3E",X"AA",X"E5",
		X"77",X"3C",X"3C",X"2B",X"77",X"2B",X"36",X"BC",X"2B",X"3E",X"B4",X"77",X"3C",X"3C",X"19",X"77",
		X"E1",X"19",X"3E",X"AF",X"77",X"3C",X"19",X"77",X"2B",X"3E",X"B8",X"77",X"3D",X"A7",X"ED",X"52",
		X"77",X"2B",X"19",X"E5",X"36",X"BE",X"19",X"3E",X"B2",X"77",X"3C",X"19",X"77",X"E1",X"2B",X"3E",
		X"A4",X"CD",X"07",X"27",X"E5",X"23",X"36",X"BD",X"19",X"3E",X"A7",X"CD",X"07",X"27",X"E1",X"3E",
		X"A4",X"CD",X"07",X"27",X"21",X"4E",X"D3",X"36",X"BF",X"2B",X"36",X"AD",X"A7",X"ED",X"52",X"36",
		X"AE",X"2B",X"3E",X"BB",X"CD",X"11",X"27",X"21",X"50",X"D3",X"36",X"93",X"23",X"36",X"F1",X"19",
		X"36",X"67",X"2B",X"36",X"61",X"C9",X"F5",X"E5",X"77",X"3C",X"E5",X"19",X"77",X"E1",X"2B",X"3C",
		X"77",X"19",X"3C",X"77",X"E1",X"F1",X"C9",X"C5",X"06",X"03",X"77",X"3C",X"19",X"10",X"FB",X"C1",
		X"C9",X"C5",X"06",X"03",X"77",X"3D",X"A7",X"ED",X"52",X"10",X"F9",X"C1",X"C9",X"06",X"09",X"21",
		X"8B",X"D1",X"DD",X"21",X"F1",X"2E",X"0E",X"03",X"CD",X"B3",X"27",X"06",X"02",X"21",X"EA",X"D1",
		X"DD",X"21",X"FA",X"2E",X"0E",X"03",X"CD",X"B3",X"27",X"06",X"0E",X"21",X"29",X"D1",X"DD",X"21",
		X"FC",X"2E",X"0E",X"07",X"CD",X"B3",X"27",X"06",X"05",X"21",X"C7",X"D1",X"DD",X"21",X"0A",X"2F",
		X"0E",X"01",X"CD",X"B3",X"27",X"3A",X"02",X"90",X"CB",X"77",X"20",X"33",X"06",X"03",X"21",X"05",
		X"D1",X"DD",X"21",X"21",X"2F",X"0E",X"01",X"CD",X"B3",X"27",X"06",X"0E",X"21",X"85",X"D1",X"DD",
		X"21",X"24",X"2F",X"CD",X"B3",X"27",X"11",X"00",X"04",X"21",X"C5",X"D0",X"0E",X"04",X"E5",X"19",
		X"71",X"E1",X"36",X"01",X"21",X"65",X"D1",X"E5",X"19",X"71",X"E1",X"36",X"02",X"18",X"23",X"3A",
		X"5E",X"60",X"FE",X"01",X"20",X"C6",X"11",X"00",X"04",X"21",X"C5",X"D0",X"0E",X"04",X"E5",X"19",
		X"71",X"E1",X"36",X"01",X"06",X"12",X"21",X"05",X"D1",X"DD",X"21",X"0F",X"2F",X"0E",X"01",X"CD",
		X"B3",X"27",X"C9",X"D5",X"11",X"00",X"04",X"E5",X"19",X"71",X"E1",X"DD",X"7E",X"00",X"77",X"D5",
		X"11",X"20",X"00",X"19",X"DD",X"23",X"D1",X"10",X"EE",X"D1",X"C9",X"F5",X"C5",X"D5",X"E5",X"06",
		X"09",X"21",X"82",X"D4",X"3E",X"02",X"11",X"20",X"00",X"77",X"23",X"77",X"19",X"77",X"2B",X"77",
		X"19",X"10",X"F6",X"18",X"07",X"F5",X"C5",X"D5",X"E5",X"11",X"20",X"00",X"3A",X"5E",X"60",X"47",
		X"3E",X"09",X"B8",X"38",X"1C",X"AF",X"21",X"03",X"90",X"ED",X"6F",X"21",X"82",X"D0",X"FE",X"0F",
		X"20",X"0B",X"0E",X"E9",X"79",X"CD",X"16",X"28",X"19",X"10",X"F9",X"18",X"04",X"0E",X"ED",X"18",
		X"F3",X"E1",X"D1",X"C1",X"F1",X"C9",X"D5",X"11",X"20",X"00",X"77",X"3D",X"23",X"77",X"3D",X"19",
		X"77",X"3D",X"2B",X"77",X"D1",X"C9",X"11",X"20",X"00",X"06",X"08",X"21",X"81",X"D6",X"3E",X"02",
		X"77",X"19",X"10",X"FC",X"3A",X"02",X"90",X"CB",X"77",X"28",X"1B",X"06",X"06",X"DD",X"21",X"81",
		X"D2",X"21",X"E7",X"2E",X"CD",X"CF",X"29",X"21",X"61",X"D3",X"3A",X"5E",X"60",X"FE",X"09",X"38",
		X"02",X"3E",X"09",X"77",X"18",X"0C",X"06",X"04",X"DD",X"21",X"01",X"D3",X"21",X"ED",X"2E",X"CD",
		X"CF",X"29",X"C9",X"F5",X"21",X"D1",X"D0",X"DD",X"21",X"32",X"2F",X"FE",X"01",X"30",X"0D",X"CD",
		X"F5",X"28",X"11",X"5E",X"00",X"19",X"DD",X"7E",X"00",X"77",X"18",X"04",X"DD",X"23",X"18",X"EF",
		X"F1",X"21",X"8F",X"D1",X"DD",X"21",X"36",X"2F",X"FE",X"01",X"F5",X"30",X"20",X"CD",X"F5",X"28",
		X"11",X"1D",X"00",X"19",X"CD",X"F5",X"28",X"11",X"23",X"00",X"19",X"CD",X"F5",X"28",X"23",X"23",
		X"CD",X"F5",X"28",X"11",X"3E",X"00",X"19",X"DD",X"7E",X"00",X"77",X"18",X"04",X"DD",X"23",X"18",
		X"DC",X"F1",X"21",X"71",X"D2",X"DD",X"21",X"40",X"2F",X"FE",X"01",X"F5",X"30",X"0D",X"CD",X"F5",
		X"28",X"11",X"3E",X"00",X"19",X"DD",X"7E",X"00",X"77",X"18",X"04",X"DD",X"23",X"18",X"EF",X"F1",
		X"21",X"EC",X"D2",X"DD",X"21",X"44",X"2F",X"FE",X"01",X"F5",X"30",X"13",X"CD",X"F5",X"28",X"23",
		X"23",X"23",X"CD",X"F5",X"28",X"11",X"40",X"00",X"19",X"DD",X"7E",X"00",X"77",X"18",X"04",X"DD",
		X"23",X"18",X"E9",X"F1",X"C9",X"DD",X"7E",X"00",X"77",X"DD",X"23",X"DD",X"23",X"C9",X"E5",X"CD",
		X"1C",X"29",X"CD",X"C1",X"2A",X"21",X"B8",X"D1",X"CD",X"E3",X"1E",X"CD",X"82",X"29",X"CD",X"A8",
		X"29",X"CD",X"DE",X"29",X"CD",X"48",X"2A",X"CD",X"A6",X"2A",X"E1",X"C9",X"21",X"B8",X"D5",X"3E",
		X"05",X"06",X"06",X"CD",X"74",X"29",X"21",X"D5",X"D5",X"3E",X"01",X"05",X"CD",X"74",X"29",X"21",
		X"74",X"D5",X"3E",X"04",X"06",X"0A",X"CD",X"74",X"29",X"21",X"33",X"D5",X"3E",X"06",X"06",X"0F",
		X"CD",X"74",X"29",X"21",X"50",X"D5",X"3E",X"06",X"06",X"0C",X"CD",X"74",X"29",X"23",X"CD",X"74",
		X"29",X"21",X"AD",X"D5",X"3E",X"05",X"06",X"06",X"CD",X"74",X"29",X"23",X"CD",X"74",X"29",X"21",
		X"AA",X"D5",X"CD",X"74",X"29",X"23",X"CD",X"74",X"29",X"21",X"88",X"D5",X"3E",X"07",X"06",X"09",
		X"CD",X"74",X"29",X"C9",X"C5",X"E5",X"F5",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"F1",X"E1",
		X"C1",X"C9",X"21",X"D5",X"D1",X"36",X"2A",X"11",X"20",X"00",X"19",X"CD",X"44",X"1F",X"DD",X"21",
		X"21",X"60",X"DD",X"36",X"00",X"82",X"DD",X"36",X"01",X"40",X"DD",X"36",X"02",X"AE",X"CD",X"7F",
		X"1F",X"DD",X"77",X"03",X"DD",X"70",X"04",X"C9",X"CD",X"26",X"1F",X"06",X"11",X"21",X"4A",X"2F",
		X"11",X"0F",X"00",X"3D",X"28",X"03",X"19",X"10",X"FA",X"DD",X"21",X"33",X"D1",X"06",X"0F",X"CD",
		X"CF",X"29",X"06",X"09",X"DD",X"21",X"88",X"D1",X"21",X"58",X"30",X"CD",X"CF",X"29",X"C9",X"D5",
		X"11",X"20",X"00",X"7E",X"DD",X"77",X"00",X"23",X"DD",X"19",X"10",X"F7",X"D1",X"C9",X"CD",X"26",
		X"1F",X"21",X"B0",X"D2",X"FE",X"12",X"38",X"07",X"06",X"06",X"CD",X"32",X"2A",X"18",X"42",X"FE",
		X"0A",X"38",X"0D",X"06",X"05",X"11",X"20",X"00",X"A7",X"ED",X"52",X"CD",X"32",X"2A",X"18",X"31",
		X"FE",X"05",X"38",X"0D",X"06",X"04",X"11",X"40",X"00",X"A7",X"ED",X"52",X"CD",X"32",X"2A",X"18",
		X"20",X"FE",X"02",X"38",X"0D",X"06",X"03",X"11",X"60",X"00",X"A7",X"ED",X"52",X"CD",X"32",X"2A",
		X"18",X"0F",X"FE",X"01",X"38",X"0B",X"06",X"02",X"11",X"80",X"00",X"A7",X"ED",X"52",X"CD",X"32",
		X"2A",X"C9",X"11",X"20",X"00",X"36",X"63",X"23",X"36",X"73",X"A7",X"ED",X"52",X"36",X"F0",X"2B",
		X"36",X"A3",X"A7",X"ED",X"52",X"10",X"EE",X"C9",X"21",X"4D",X"D2",X"FD",X"21",X"6F",X"60",X"06",
		X"03",X"DD",X"21",X"AD",X"0C",X"FD",X"23",X"FD",X"5E",X"00",X"CB",X"23",X"CB",X"23",X"16",X"00",
		X"DD",X"19",X"CD",X"68",X"2A",X"10",X"EA",X"C9",X"D5",X"11",X"20",X"00",X"DD",X"7E",X"00",X"77",
		X"23",X"DD",X"23",X"DD",X"7E",X"00",X"3C",X"77",X"A7",X"ED",X"52",X"CD",X"91",X"2A",X"77",X"2B",
		X"DD",X"23",X"DD",X"23",X"DD",X"7E",X"00",X"3C",X"77",X"11",X"20",X"00",X"A7",X"ED",X"52",X"D1",
		X"C9",X"C5",X"FD",X"7E",X"00",X"06",X"F1",X"FE",X"09",X"28",X"08",X"D6",X"05",X"38",X"04",X"3C",
		X"80",X"18",X"01",X"78",X"C1",X"C9",X"21",X"4A",X"D2",X"06",X"03",X"11",X"20",X"00",X"36",X"62",
		X"23",X"36",X"71",X"A7",X"ED",X"52",X"36",X"EF",X"2B",X"36",X"A1",X"A7",X"ED",X"52",X"10",X"EE",
		X"C9",X"06",X"15",X"21",X"A6",X"D0",X"3E",X"32",X"77",X"CD",X"FB",X"2A",X"23",X"10",X"F9",X"36",
		X"30",X"CD",X"FB",X"2A",X"06",X"15",X"21",X"DB",X"D0",X"11",X"20",X"00",X"3D",X"77",X"CD",X"FB",
		X"2A",X"19",X"10",X"F9",X"21",X"C6",X"D0",X"11",X"20",X"00",X"3E",X"FF",X"0E",X"15",X"E5",X"06",
		X"15",X"77",X"19",X"10",X"FC",X"E1",X"23",X"0D",X"20",X"F4",X"C9",X"E5",X"D5",X"11",X"00",X"04",
		X"19",X"36",X"00",X"D1",X"E1",X"C9",X"01",X"FF",X"03",X"21",X"00",X"D4",X"AF",X"77",X"23",X"0B",
		X"78",X"B1",X"20",X"F8",X"C9",X"3A",X"65",X"60",X"FE",X"00",X"20",X"06",X"DD",X"21",X"A3",X"60",
		X"18",X"04",X"DD",X"21",X"A6",X"60",X"3E",X"01",X"DD",X"4E",X"00",X"DD",X"56",X"01",X"DD",X"5E",
		X"02",X"06",X"00",X"CB",X"3B",X"CB",X"1A",X"CB",X"19",X"CB",X"10",X"CD",X"6E",X"2B",X"F5",X"FE",
		X"03",X"28",X"1C",X"FE",X"05",X"28",X"18",X"FE",X"06",X"28",X"14",X"FE",X"0A",X"28",X"10",X"FE",
		X"0C",X"28",X"0C",X"FE",X"0D",X"28",X"08",X"FE",X"0F",X"28",X"04",X"FE",X"10",X"20",X"04",X"CB",
		X"18",X"CB",X"15",X"F1",X"3C",X"FE",X"15",X"20",X"C8",X"4D",X"CD",X"1C",X"2C",X"C9",X"D5",X"C5",
		X"DD",X"E5",X"F5",X"E5",X"5F",X"4F",X"CD",X"04",X"2C",X"78",X"FE",X"00",X"20",X"1A",X"36",X"36",
		X"E5",X"23",X"36",X"39",X"E1",X"2B",X"36",X"FF",X"11",X"20",X"00",X"23",X"E5",X"19",X"36",X"37",
		X"E1",X"A7",X"ED",X"52",X"36",X"35",X"18",X"18",X"36",X"3E",X"E5",X"23",X"36",X"3D",X"E1",X"2B",
		X"36",X"3F",X"11",X"20",X"00",X"23",X"E5",X"19",X"36",X"FF",X"E1",X"A7",X"ED",X"52",X"36",X"40",
		X"19",X"E5",X"FD",X"21",X"45",X"0D",X"DD",X"21",X"55",X"0D",X"16",X"00",X"59",X"1D",X"D5",X"CB",
		X"3B",X"DD",X"19",X"DD",X"4E",X"00",X"D1",X"CB",X"43",X"20",X"06",X"79",X"E6",X"0F",X"4F",X"18",
		X"08",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"CB",X"39",X"C5",X"06",X"00",X"CB",X"21",X"CB",X"21",
		X"FD",X"09",X"C1",X"78",X"FE",X"00",X"20",X"04",X"FD",X"23",X"FD",X"23",X"01",X"40",X"00",X"A7",
		X"ED",X"42",X"FD",X"7E",X"00",X"77",X"E1",X"23",X"23",X"FD",X"7E",X"01",X"77",X"E1",X"F1",X"DD",
		X"E1",X"C1",X"D1",X"C9",X"D5",X"DD",X"E5",X"DD",X"21",X"1D",X"0D",X"16",X"00",X"1D",X"CB",X"23",
		X"DD",X"19",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"DD",X"E1",X"D1",X"C9",X"16",X"00",X"CB",X"21",
		X"CB",X"12",X"CB",X"21",X"CB",X"12",X"21",X"2F",X"D1",X"CD",X"5A",X"2C",X"CB",X"21",X"CB",X"12",
		X"CB",X"21",X"CB",X"12",X"21",X"77",X"D1",X"CD",X"5A",X"2C",X"1E",X"00",X"CB",X"21",X"CB",X"12",
		X"CB",X"21",X"CB",X"13",X"CB",X"21",X"CB",X"12",X"CB",X"21",X"CB",X"13",X"21",X"6F",X"D2",X"CD",
		X"5A",X"2C",X"53",X"21",X"75",X"D2",X"CD",X"5A",X"2C",X"C9",X"7A",X"FE",X"00",X"28",X"0C",X"FE",
		X"02",X"28",X"0C",X"FE",X"03",X"20",X"0A",X"36",X"3B",X"18",X"06",X"36",X"34",X"18",X"02",X"36",
		X"3A",X"16",X"00",X"C9",X"CD",X"C1",X"2A",X"21",X"26",X"60",X"CB",X"4E",X"28",X"03",X"CD",X"A2",
		X"2C",X"21",X"50",X"D1",X"3E",X"FF",X"06",X"0D",X"CD",X"7D",X"1E",X"21",X"50",X"D5",X"3E",X"06",
		X"06",X"0D",X"CD",X"7D",X"1E",X"21",X"6D",X"0D",X"DD",X"21",X"50",X"D1",X"06",X"0D",X"CD",X"CF",
		X"29",X"C9",X"AF",X"21",X"21",X"60",X"77",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"21",X"2B",X"60",
		X"06",X"07",X"11",X"05",X"00",X"AF",X"77",X"D5",X"CD",X"4F",X"2E",X"D1",X"19",X"10",X"F7",X"21",
		X"26",X"60",X"E5",X"36",X"12",X"23",X"CD",X"4F",X"2E",X"35",X"7E",X"FE",X"07",X"20",X"F7",X"E1",
		X"36",X"22",X"23",X"23",X"CD",X"4F",X"2E",X"35",X"7E",X"FE",X"22",X"20",X"F7",X"21",X"26",X"60",
		X"36",X"00",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"3A",X"65",X"60",X"FE",X"00",X"28",X"05",X"21",
		X"67",X"60",X"18",X"03",X"21",X"66",X"60",X"34",X"CD",X"77",X"1D",X"C9",X"F5",X"CD",X"C1",X"2A",
		X"21",X"71",X"D5",X"06",X"0A",X"3E",X"07",X"CD",X"7D",X"1E",X"2B",X"CD",X"7D",X"1E",X"2B",X"CD",
		X"7D",X"1E",X"F1",X"FE",X"01",X"28",X"10",X"30",X"28",X"06",X"09",X"DD",X"21",X"90",X"D1",X"21",
		X"68",X"0E",X"CD",X"CF",X"29",X"18",X"32",X"06",X"0A",X"DD",X"21",X"71",X"D1",X"21",X"71",X"0E",
		X"CD",X"CF",X"29",X"06",X"09",X"DD",X"21",X"8F",X"D1",X"21",X"68",X"0E",X"CD",X"CF",X"29",X"18",
		X"18",X"06",X"0A",X"DD",X"21",X"71",X"D1",X"21",X"7B",X"0E",X"CD",X"CF",X"29",X"06",X"09",X"DD",
		X"21",X"8F",X"D1",X"21",X"68",X"0E",X"CD",X"CF",X"29",X"C9",X"F5",X"3A",X"02",X"90",X"CB",X"67",
		X"28",X"F9",X"F1",X"C9",X"21",X"26",X"60",X"36",X"82",X"06",X"1E",X"3E",X"E4",X"23",X"23",X"23",
		X"CD",X"4F",X"2E",X"77",X"23",X"36",X"00",X"2B",X"10",X"F6",X"06",X"06",X"C6",X"04",X"0E",X"05",
		X"77",X"CD",X"4F",X"2E",X"0D",X"20",X"F9",X"10",X"F3",X"06",X"06",X"3E",X"48",X"0E",X"05",X"77",
		X"23",X"36",X"09",X"CB",X"E6",X"2B",X"CD",X"4F",X"2E",X"0D",X"20",X"F3",X"C6",X"04",X"10",X"ED",
		X"06",X"1E",X"77",X"CD",X"4F",X"2E",X"10",X"FA",X"DD",X"21",X"02",X"60",X"DD",X"CB",X"00",X"C6",
		X"2B",X"11",X"CE",X"2D",X"D5",X"CD",X"D7",X"2D",X"CD",X"14",X"2E",X"CD",X"14",X"2E",X"CD",X"D7",
		X"2D",X"CD",X"D7",X"2D",X"CD",X"14",X"2E",X"CD",X"14",X"2E",X"CD",X"D7",X"2D",X"D1",X"21",X"26",
		X"60",X"36",X"00",X"CD",X"2F",X"3F",X"C9",X"2B",X"06",X"02",X"3E",X"AF",X"34",X"BE",X"CA",X"12",
		X"2E",X"CD",X"4F",X"2E",X"10",X"F6",X"06",X"04",X"3E",X"AF",X"34",X"BE",X"CA",X"12",X"2E",X"23",
		X"34",X"3E",X"D7",X"BE",X"CA",X"12",X"2E",X"CD",X"4F",X"2E",X"2B",X"10",X"EB",X"23",X"06",X"04",
		X"34",X"BE",X"CA",X"12",X"2E",X"CD",X"4F",X"2E",X"10",X"F6",X"06",X"05",X"CD",X"4F",X"2E",X"10",
		X"FB",X"C9",X"D1",X"C9",X"2B",X"06",X"02",X"AF",X"35",X"BE",X"CA",X"4D",X"2E",X"CD",X"4F",X"2E",
		X"10",X"F6",X"06",X"04",X"AF",X"35",X"BE",X"CA",X"4D",X"2E",X"23",X"34",X"3E",X"D7",X"BE",X"CA",
		X"4D",X"2E",X"CD",X"4F",X"2E",X"2B",X"10",X"EC",X"23",X"06",X"04",X"34",X"BE",X"CA",X"4D",X"2E",
		X"CD",X"4F",X"2E",X"10",X"F6",X"06",X"05",X"CD",X"4F",X"2E",X"10",X"FB",X"C9",X"D1",X"C9",X"F5",
		X"E5",X"C5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"C1",X"E1",X"F1",X"C9",X"21",X"A4",X"0E",X"CD",
		X"26",X"1F",X"CB",X"47",X"20",X"01",X"23",X"3A",X"B9",X"61",X"BE",X"DA",X"9E",X"2E",X"3A",X"65",
		X"60",X"FE",X"00",X"28",X"0C",X"3A",X"02",X"90",X"CB",X"6F",X"28",X"05",X"3A",X"01",X"90",X"18",
		X"03",X"3A",X"00",X"90",X"FE",X"00",X"CA",X"9E",X"2E",X"3A",X"98",X"61",X"21",X"C4",X"61",X"06",
		X"04",X"CB",X"3F",X"30",X"02",X"CB",X"DF",X"77",X"23",X"10",X"F6",X"C3",X"CB",X"2E",X"21",X"C4",
		X"61",X"06",X"04",X"ED",X"5F",X"E6",X"0F",X"CB",X"3F",X"3C",X"FE",X"03",X"38",X"0D",X"FE",X"05",
		X"38",X"0E",X"FE",X"07",X"38",X"0F",X"3E",X"08",X"C3",X"C7",X"2E",X"3E",X"01",X"C3",X"C7",X"2E",
		X"3E",X"02",X"C3",X"C7",X"2E",X"3E",X"04",X"77",X"23",X"10",X"D8",X"CD",X"D8",X"46",X"C9",X"18",
		X"19",X"17",X"0D",X"1B",X"0D",X"1D",X"11",X"1D",X"18",X"0D",X"0A",X"22",X"2E",X"1C",X"FF",X"11",
		X"12",X"FF",X"1C",X"0C",X"18",X"1B",X"0E",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"0F",X"1B",X"0E",
		X"0E",X"19",X"1B",X"0E",X"1C",X"0E",X"17",X"1D",X"0E",X"0D",X"0B",X"22",X"1E",X"17",X"12",X"1F",
		X"0E",X"1B",X"1C",X"0A",X"15",X"2F",X"01",X"09",X"08",X"01",X"19",X"1B",X"0E",X"1C",X"1C",X"19",
		X"15",X"0A",X"22",X"0E",X"1B",X"FF",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"FF",X"18",X"17",X"15",
		X"22",X"18",X"1B",X"FF",X"FF",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"FF",X"0B",X"1E",X"1D",X"1D",
		X"18",X"17",X"C0",X"AB",X"C1",X"A8",X"A8",X"C1",X"B9",X"C3",X"B2",X"C2",X"AB",X"C0",X"BD",X"C4",
		X"C5",X"AF",X"C2",X"B2",X"B9",X"C3",X"BD",X"C4",X"A8",X"C1",X"FF",X"FF",X"FF",X"0C",X"1E",X"0C",
		X"1E",X"16",X"0B",X"0E",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0E",X"10",X"10",X"FF",
		X"19",X"15",X"0A",X"17",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"0A",X"1B",X"1B",
		X"18",X"1D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1B",X"0A",X"0D",X"12",X"1C",
		X"11",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"19",X"0A",X"1B",X"1C",X"15",X"0E",
		X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1D",X"18",X"16",X"0A",X"1D",X"18",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"19",X"1E",X"16",X"19",X"14",X"12",X"17",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0B",X"0A",X"16",X"0B",X"18",X"18",X"FF",X"1C",X"11",X"18",X"18",X"1D",
		X"FF",X"FF",X"13",X"0A",X"19",X"0A",X"17",X"0E",X"1C",X"0E",X"FF",X"1B",X"0A",X"0D",X"12",X"1C",
		X"11",X"FF",X"FF",X"FF",X"16",X"1E",X"1C",X"11",X"1B",X"18",X"18",X"16",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"19",X"18",X"1D",X"0A",X"1D",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"18",X"17",X"12",X"18",X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",X"11",
		X"12",X"17",X"0E",X"1C",X"0E",X"FF",X"0C",X"0A",X"0B",X"0B",X"0A",X"10",X"0E",X"FF",X"FF",X"FF",
		X"FF",X"1D",X"1E",X"1B",X"17",X"12",X"19",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1B",
		X"0E",X"0D",X"FF",X"19",X"0E",X"19",X"0E",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0C",
		X"0E",X"15",X"0E",X"1B",X"22",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1C",X"20",X"0E",X"0E",X"1D",
		X"FF",X"19",X"18",X"1D",X"0A",X"1D",X"18",X"FF",X"FF",X"FF",X"FF",X"11",X"18",X"1B",X"1C",X"0E",
		X"1B",X"0A",X"0D",X"12",X"1C",X"11",X"FF",X"FF",X"10",X"18",X"18",X"0D",X"FF",X"15",X"1E",X"0C",
		X"14",X"79",X"DD",X"21",X"2B",X"60",X"CB",X"27",X"CB",X"27",X"81",X"16",X"00",X"5F",X"DD",X"19",
		X"DD",X"36",X"00",X"82",X"DD",X"36",X"01",X"58",X"DD",X"36",X"02",X"86",X"79",X"CD",X"87",X"30",
		X"DD",X"77",X"03",X"DD",X"70",X"04",X"C9",X"F5",X"CD",X"26",X"1F",X"FE",X"09",X"30",X"20",X"4F",
		X"FE",X"03",X"28",X"06",X"FE",X"04",X"28",X"05",X"18",X"04",X"3C",X"18",X"01",X"3D",X"47",X"79",
		X"3D",X"E5",X"21",X"8B",X"0C",X"16",X"00",X"5F",X"19",X"7E",X"4F",X"E1",X"F1",X"79",X"C9",X"3D",
		X"E6",X"07",X"FE",X"05",X"38",X"02",X"D6",X"05",X"47",X"F1",X"80",X"47",X"04",X"4F",X"3E",X"18",
		X"CB",X"21",X"CB",X"21",X"CB",X"21",X"08",X"79",X"CB",X"21",X"81",X"4F",X"08",X"81",X"C9",X"CD",
		X"A9",X"34",X"47",X"3E",X"75",X"90",X"32",X"A9",X"60",X"C9",X"06",X"03",X"3A",X"65",X"60",X"FE",
		X"00",X"28",X"05",X"21",X"A6",X"60",X"18",X"03",X"21",X"A3",X"60",X"36",X"95",X"23",X"36",X"6A",
		X"23",X"36",X"0A",X"C9",X"3A",X"65",X"60",X"FE",X"00",X"28",X"05",X"3A",X"A0",X"60",X"18",X"03",
		X"3A",X"9D",X"60",X"06",X"07",X"21",X"BD",X"D4",X"16",X"03",X"1E",X"07",X"1F",X"38",X"03",X"73",
		X"18",X"01",X"72",X"D5",X"11",X"20",X"00",X"19",X"D1",X"10",X"F1",X"C9",X"3A",X"65",X"60",X"FE",
		X"00",X"28",X"05",X"3A",X"A1",X"60",X"18",X"03",X"3A",X"9E",X"60",X"06",X"05",X"21",X"DD",X"D5",
		X"16",X"03",X"1E",X"06",X"1F",X"38",X"03",X"73",X"18",X"01",X"72",X"D5",X"11",X"20",X"00",X"19",
		X"D1",X"10",X"F1",X"C9",X"21",X"9F",X"60",X"3A",X"65",X"60",X"FE",X"00",X"28",X"03",X"21",X"A2",
		X"60",X"AF",X"77",X"C9",X"3A",X"65",X"60",X"FE",X"00",X"28",X"05",X"3A",X"A2",X"60",X"18",X"03",
		X"3A",X"9F",X"60",X"21",X"BD",X"D6",X"11",X"20",X"00",X"06",X"03",X"0E",X"05",X"FE",X"00",X"20",
		X"0D",X"70",X"19",X"70",X"19",X"70",X"19",X"70",X"19",X"70",X"19",X"70",X"18",X"13",X"71",X"19",
		X"71",X"FE",X"01",X"28",X"EF",X"19",X"71",X"19",X"71",X"FE",X"02",X"28",X"EB",X"19",X"71",X"19",
		X"71",X"C9",X"CD",X"63",X"33",X"CD",X"3D",X"3F",X"06",X"0A",X"16",X"00",X"FD",X"21",X"91",X"60",
		X"FD",X"E5",X"FD",X"7E",X"01",X"CD",X"C5",X"32",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",
		X"14",X"3E",X"03",X"BA",X"20",X"EC",X"CD",X"A9",X"34",X"FD",X"E1",X"06",X"0B",X"16",X"00",X"08",
		X"FD",X"7E",X"02",X"CD",X"C5",X"32",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"14",X"08",
		X"3D",X"28",X"0E",X"08",X"7A",X"FE",X"03",X"20",X"E7",X"FD",X"21",X"92",X"60",X"16",X"00",X"18",
		X"DF",X"16",X"00",X"FD",X"21",X"70",X"60",X"ED",X"5F",X"07",X"CB",X"12",X"07",X"E6",X"03",X"8A",
		X"16",X"00",X"FE",X"01",X"28",X"32",X"38",X"10",X"FE",X"03",X"CA",X"68",X"32",X"DA",X"48",X"32",
		X"FE",X"05",X"CA",X"A7",X"32",X"C3",X"88",X"32",X"FD",X"46",X"00",X"3A",X"91",X"60",X"CD",X"C5",
		X"32",X"14",X"FD",X"46",X"01",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"02",X"3A",
		X"99",X"60",X"CD",X"C5",X"32",X"C3",X"C4",X"32",X"FD",X"46",X"00",X"3A",X"91",X"60",X"CD",X"C5",
		X"32",X"14",X"FD",X"46",X"02",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"01",X"3A",
		X"99",X"60",X"CD",X"C5",X"32",X"C3",X"C4",X"32",X"FD",X"46",X"01",X"3A",X"91",X"60",X"CD",X"C5",
		X"32",X"14",X"FD",X"46",X"00",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"02",X"3A",
		X"99",X"60",X"CD",X"C5",X"32",X"C3",X"C4",X"32",X"FD",X"46",X"01",X"3A",X"91",X"60",X"CD",X"C5",
		X"32",X"14",X"FD",X"46",X"02",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"00",X"3A",
		X"99",X"60",X"CD",X"C5",X"32",X"C3",X"C4",X"32",X"FD",X"46",X"02",X"3A",X"91",X"60",X"CD",X"C5",
		X"32",X"14",X"FD",X"46",X"00",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"01",X"3A",
		X"99",X"60",X"CD",X"C5",X"32",X"18",X"1D",X"FD",X"46",X"02",X"3A",X"91",X"60",X"CD",X"C5",X"32",
		X"14",X"FD",X"46",X"01",X"3A",X"95",X"60",X"CD",X"C5",X"32",X"14",X"FD",X"46",X"00",X"3A",X"99",
		X"60",X"CD",X"C5",X"32",X"C9",X"F5",X"CD",X"79",X"3A",X"CD",X"44",X"34",X"F1",X"F5",X"C5",X"4F",
		X"7A",X"CD",X"3B",X"33",X"C1",X"78",X"18",X"01",X"F5",X"C5",X"06",X"07",X"FE",X"0A",X"20",X"06",
		X"DD",X"21",X"A5",X"0C",X"18",X"0A",X"FE",X"0B",X"20",X"09",X"06",X"06",X"DD",X"21",X"A9",X"0C",
		X"D5",X"18",X"0E",X"DD",X"21",X"AD",X"0C",X"D5",X"CB",X"27",X"CB",X"27",X"16",X"00",X"5F",X"DD",
		X"19",X"DD",X"7E",X"00",X"77",X"11",X"00",X"04",X"E5",X"19",X"70",X"E1",X"DD",X"7E",X"01",X"23",
		X"CB",X"49",X"28",X"01",X"3C",X"77",X"E5",X"19",X"70",X"E1",X"D5",X"11",X"E0",X"FF",X"19",X"D1",
		X"DD",X"7E",X"02",X"81",X"77",X"E5",X"19",X"70",X"E1",X"2B",X"DD",X"7E",X"03",X"CB",X"41",X"28",
		X"01",X"3C",X"77",X"E5",X"19",X"70",X"E1",X"D1",X"C1",X"F1",X"C9",X"DD",X"E5",X"C5",X"FE",X"01",
		X"28",X"0C",X"38",X"05",X"21",X"34",X"0C",X"18",X"08",X"21",X"02",X"0C",X"18",X"03",X"21",X"16",
		X"0C",X"06",X"00",X"CB",X"21",X"09",X"E5",X"DD",X"E1",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"C1",
		X"DD",X"E1",X"C9",X"06",X"04",X"21",X"91",X"60",X"E5",X"DD",X"E1",X"ED",X"5F",X"4F",X"E6",X"07",
		X"CB",X"21",X"CE",X"00",X"CB",X"21",X"CE",X"00",X"CD",X"A2",X"33",X"38",X"EE",X"77",X"23",X"10",
		X"EA",X"21",X"95",X"60",X"06",X"02",X"C5",X"E5",X"DD",X"E1",X"06",X"04",X"ED",X"5F",X"4F",X"E6",
		X"0F",X"FE",X"0F",X"28",X"F7",X"CD",X"A2",X"33",X"38",X"F2",X"77",X"23",X"10",X"EE",X"C1",X"10",
		X"E5",X"C9",X"08",X"78",X"FE",X"01",X"20",X"14",X"08",X"DD",X"BE",X"02",X"28",X"1F",X"DD",X"BE",
		X"01",X"28",X"1A",X"DD",X"BE",X"00",X"28",X"15",X"37",X"3F",X"18",X"12",X"FE",X"02",X"20",X"03",
		X"08",X"18",X"EB",X"FE",X"03",X"20",X"03",X"08",X"18",X"E9",X"08",X"18",X"EB",X"37",X"C9",X"DD",
		X"21",X"6E",X"60",X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"DD",X"34",X"00",X"18",X"03",X"DD",
		X"34",X"01",X"C9",X"21",X"C6",X"D0",X"CD",X"25",X"34",X"D5",X"11",X"06",X"00",X"19",X"D1",X"E5",
		X"DD",X"E1",X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"06",X"DD",X"77",X"08",X"DD",X"77",
		X"0A",X"DD",X"77",X"0C",X"DD",X"77",X"0E",X"DD",X"19",X"DD",X"71",X"00",X"DD",X"71",X"02",X"DD",
		X"71",X"06",X"DD",X"71",X"08",X"DD",X"71",X"0A",X"DD",X"71",X"0C",X"DD",X"71",X"0E",X"21",X"46",
		X"D2",X"CD",X"25",X"34",X"C9",X"0E",X"02",X"3E",X"E5",X"11",X"00",X"04",X"06",X"05",X"C5",X"06",
		X"0B",X"77",X"E5",X"19",X"71",X"E1",X"23",X"23",X"10",X"F7",X"D5",X"11",X"2A",X"00",X"19",X"D1",
		X"C1",X"10",X"EB",X"C9",X"0E",X"00",X"FE",X"0A",X"28",X"5E",X"FE",X"64",X"28",X"5A",X"FE",X"07",
		X"38",X"24",X"FE",X"09",X"28",X"20",X"FE",X"31",X"28",X"1C",X"FE",X"3A",X"28",X"18",X"FE",X"3C",
		X"28",X"14",X"FE",X"43",X"28",X"10",X"FE",X"5A",X"28",X"0C",X"FE",X"6B",X"28",X"08",X"FE",X"6D",
		X"28",X"04",X"FE",X"6E",X"20",X"03",X"0C",X"18",X"2E",X"FE",X"18",X"28",X"28",X"FE",X"1C",X"28",
		X"24",X"FE",X"2C",X"28",X"20",X"FE",X"3A",X"28",X"1C",X"FE",X"3B",X"28",X"18",X"FE",X"3E",X"28",
		X"14",X"FE",X"56",X"28",X"10",X"FE",X"6A",X"28",X"0C",X"FE",X"6C",X"28",X"08",X"FE",X"6F",X"28",
		X"04",X"FE",X"70",X"20",X"02",X"0C",X"0C",X"0C",X"C9",X"CD",X"26",X"1F",X"FE",X"01",X"20",X"04",
		X"3E",X"02",X"18",X"1A",X"FE",X"05",X"30",X"04",X"3E",X"03",X"18",X"12",X"FE",X"0A",X"30",X"04",
		X"3E",X"04",X"18",X"0A",X"FE",X"11",X"30",X"04",X"3E",X"05",X"18",X"02",X"3E",X"06",X"C9",X"C5",
		X"E5",X"FD",X"7E",X"00",X"FE",X"0C",X"38",X"1B",X"FE",X"FF",X"28",X"06",X"FE",X"E5",X"28",X"02",
		X"3E",X"FF",X"77",X"FE",X"FF",X"28",X"26",X"11",X"00",X"04",X"19",X"36",X"02",X"21",X"A9",X"60",
		X"34",X"18",X"1A",X"FE",X"0B",X"28",X"06",X"E5",X"21",X"A9",X"60",X"34",X"E1",X"41",X"08",X"79",
		X"CD",X"44",X"34",X"08",X"47",X"CD",X"D8",X"32",X"E1",X"E5",X"CD",X"7B",X"3F",X"E1",X"C1",X"C9",
		X"0E",X"00",X"21",X"C6",X"D0",X"3A",X"65",X"60",X"FE",X"00",X"28",X"06",X"DD",X"21",X"21",X"61",
		X"18",X"04",X"DD",X"21",X"AC",X"60",X"06",X"0B",X"CD",X"63",X"35",X"DD",X"77",X"00",X"DD",X"23",
		X"0C",X"79",X"FE",X"37",X"20",X"20",X"11",X"32",X"00",X"19",X"CD",X"63",X"35",X"DD",X"77",X"00",
		X"DD",X"23",X"0C",X"23",X"23",X"CD",X"63",X"35",X"DD",X"77",X"00",X"DD",X"23",X"0C",X"06",X"05",
		X"23",X"23",X"23",X"23",X"18",X"D2",X"FE",X"75",X"28",X"08",X"10",X"F6",X"11",X"2C",X"00",X"19",
		X"18",X"C4",X"C9",X"FD",X"21",X"5F",X"0D",X"16",X"00",X"7E",X"FD",X"BE",X"00",X"28",X"10",X"FD",
		X"23",X"14",X"18",X"F6",X"7A",X"FE",X"01",X"28",X"02",X"30",X"14",X"FD",X"7E",X"00",X"C9",X"FE",
		X"5C",X"20",X"F1",X"E5",X"23",X"7E",X"E1",X"FE",X"66",X"38",X"E9",X"14",X"14",X"18",X"E5",X"D6",
		X"02",X"C9",X"CD",X"BC",X"3F",X"AF",X"32",X"A9",X"60",X"3A",X"65",X"60",X"FE",X"00",X"20",X"06",
		X"FD",X"21",X"AC",X"60",X"18",X"04",X"FD",X"21",X"21",X"61",X"21",X"C6",X"D0",X"0E",X"00",X"06",
		X"0B",X"CD",X"CF",X"34",X"FD",X"23",X"0C",X"79",X"FE",X"37",X"20",X"1A",X"11",X"32",X"00",X"19",
		X"CD",X"CF",X"34",X"FD",X"23",X"0C",X"23",X"23",X"CD",X"CF",X"34",X"FD",X"23",X"0C",X"06",X"05",
		X"23",X"23",X"23",X"23",X"18",X"DB",X"FE",X"75",X"28",X"08",X"10",X"F6",X"11",X"2C",X"00",X"19",
		X"18",X"CD",X"C9",X"CD",X"26",X"1F",X"21",X"AA",X"60",X"FE",X"02",X"30",X"04",X"36",X"09",X"18",
		X"0A",X"FE",X"05",X"30",X"04",X"36",X"06",X"18",X"02",X"36",X"03",X"7E",X"23",X"77",X"C9",X"21",
		X"5F",X"60",X"CB",X"66",X"CA",X"29",X"36",X"2A",X"D8",X"61",X"3A",X"27",X"60",X"E6",X"0F",X"FE",
		X"08",X"20",X"13",X"3A",X"28",X"60",X"E6",X"0F",X"FE",X"06",X"20",X"0A",X"23",X"7E",X"FE",X"FF",
		X"20",X"01",X"2B",X"22",X"D8",X"61",X"7E",X"18",X"17",X"3A",X"65",X"60",X"FE",X"00",X"28",X"0C",
		X"3A",X"02",X"90",X"CB",X"6F",X"28",X"05",X"3A",X"01",X"90",X"18",X"03",X"3A",X"00",X"90",X"2F",
		X"E6",X"0F",X"C8",X"FE",X"01",X"28",X"0B",X"FE",X"02",X"28",X"07",X"FE",X"04",X"28",X"03",X"FE",
		X"08",X"C0",X"57",X"3A",X"5F",X"60",X"CB",X"7F",X"CA",X"C1",X"36",X"3A",X"27",X"60",X"E6",X"0F",
		X"FE",X"08",X"CA",X"43",X"49",X"3A",X"28",X"60",X"E6",X"0F",X"FE",X"06",X"C2",X"4B",X"49",X"D5",
		X"AF",X"32",X"E0",X"61",X"C3",X"CE",X"36",X"CB",X"3F",X"BA",X"C2",X"1E",X"38",X"21",X"27",X"60",
		X"E6",X"0A",X"28",X"1E",X"7E",X"E6",X"0F",X"FE",X"08",X"38",X"03",X"35",X"18",X"01",X"34",X"23",
		X"CB",X"5A",X"20",X"07",X"35",X"3E",X"02",X"32",X"98",X"61",X"C9",X"34",X"3E",X"08",X"32",X"98",
		X"61",X"C9",X"23",X"7E",X"E6",X"0F",X"FE",X"07",X"38",X"03",X"35",X"18",X"01",X"34",X"2B",X"CB",
		X"52",X"28",X"07",X"34",X"3E",X"04",X"32",X"98",X"61",X"C9",X"35",X"3E",X"01",X"32",X"98",X"61",
		X"C9",X"D5",X"AF",X"32",X"E0",X"61",X"3A",X"98",X"61",X"E6",X"0A",X"C2",X"6E",X"37",X"3A",X"27",
		X"60",X"47",X"3A",X"28",X"60",X"CD",X"DA",X"36",X"18",X"1B",X"D6",X"36",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"27",X"21",X"E4",X"0D",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",
		X"3E",X"08",X"0E",X"10",X"C9",X"CB",X"3A",X"CB",X"1B",X"38",X"03",X"81",X"18",X"F7",X"CD",X"03",
		X"37",X"18",X"03",X"B8",X"3F",X"C9",X"28",X"06",X"38",X"08",X"CB",X"FA",X"18",X"ED",X"67",X"6F",
		X"18",X"0D",X"67",X"CB",X"23",X"CB",X"12",X"91",X"CB",X"23",X"CB",X"12",X"30",X"F9",X"6F",X"3A",
		X"27",X"60",X"08",X"DD",X"21",X"96",X"61",X"7C",X"D6",X"04",X"57",X"08",X"BA",X"30",X"33",X"08",
		X"7A",X"D6",X"02",X"57",X"08",X"BA",X"30",X"25",X"08",X"7D",X"C6",X"05",X"5F",X"08",X"BB",X"38",
		X"17",X"08",X"7B",X"C6",X"02",X"5F",X"08",X"BB",X"D2",X"0A",X"38",X"DD",X"75",X"00",X"E5",X"21",
		X"E0",X"61",X"CB",X"CE",X"E1",X"C3",X"0A",X"38",X"DD",X"75",X"00",X"18",X"08",X"DD",X"74",X"00",
		X"18",X"EC",X"DD",X"74",X"00",X"3A",X"28",X"60",X"DD",X"77",X"01",X"C3",X"06",X"38",X"3A",X"28",
		X"60",X"47",X"3A",X"27",X"60",X"CD",X"7A",X"37",X"18",X"1B",X"D6",X"08",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"27",X"21",X"FA",X"0D",X"16",X"00",X"5F",X"19",X"5E",X"23",X"56",
		X"3E",X"36",X"0E",X"10",X"C9",X"CB",X"3A",X"CB",X"1B",X"38",X"03",X"81",X"18",X"F7",X"CD",X"03",
		X"37",X"28",X"06",X"38",X"08",X"CB",X"FA",X"18",X"F2",X"67",X"6F",X"18",X"0D",X"67",X"CB",X"23",
		X"CB",X"12",X"91",X"CB",X"23",X"CB",X"12",X"30",X"F9",X"6F",X"3A",X"28",X"60",X"08",X"DD",X"21",
		X"96",X"61",X"7C",X"D6",X"04",X"57",X"08",X"BA",X"30",X"33",X"08",X"7A",X"D6",X"03",X"57",X"08",
		X"BA",X"30",X"25",X"08",X"7D",X"C6",X"05",X"5F",X"08",X"BB",X"38",X"17",X"08",X"7B",X"C6",X"03",
		X"5F",X"08",X"BB",X"D2",X"0A",X"38",X"DD",X"75",X"01",X"E5",X"21",X"E0",X"61",X"CB",X"C6",X"E1",
		X"C3",X"0A",X"38",X"DD",X"75",X"01",X"18",X"08",X"DD",X"74",X"01",X"18",X"EC",X"DD",X"74",X"01",
		X"3A",X"27",X"60",X"DD",X"77",X"00",X"D1",X"C3",X"8C",X"38",X"D1",X"21",X"5F",X"60",X"CB",X"BE",
		X"3A",X"26",X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"BA",X"28",X"0F",X"7A",X"CB",
		X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"F6",X"02",X"32",X"26",X"60",X"C9",X"3E",X"05",X"A2",
		X"28",X"0A",X"3A",X"98",X"61",X"E6",X"05",X"CA",X"69",X"38",X"18",X"08",X"3A",X"98",X"61",X"E6",
		X"0A",X"CA",X"69",X"38",X"DD",X"21",X"27",X"60",X"7A",X"FE",X"02",X"38",X"0B",X"28",X"0E",X"FE",
		X"04",X"28",X"0F",X"DD",X"34",X"01",X"18",X"0D",X"DD",X"35",X"00",X"18",X"08",X"DD",X"35",X"01",
		X"18",X"03",X"DD",X"34",X"00",X"32",X"98",X"61",X"C9",X"3A",X"E0",X"61",X"FE",X"00",X"C8",X"CB",
		X"47",X"28",X"0D",X"21",X"28",X"60",X"3A",X"97",X"61",X"BE",X"38",X"02",X"34",X"C9",X"35",X"C9",
		X"21",X"27",X"60",X"3A",X"96",X"61",X"BE",X"38",X"F5",X"C3",X"7C",X"38",X"21",X"5F",X"60",X"CB",
		X"FE",X"3A",X"26",X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"BA",X"C2",X"1E",X"38",
		X"FD",X"21",X"26",X"60",X"DD",X"21",X"96",X"61",X"3A",X"28",X"60",X"DD",X"BE",X"01",X"20",X"36",
		X"3A",X"27",X"60",X"DD",X"BE",X"00",X"20",X"07",X"CD",X"0D",X"39",X"D2",X"44",X"38",X"C9",X"3A",
		X"27",X"60",X"DD",X"BE",X"00",X"38",X"10",X"3E",X"05",X"A2",X"C2",X"44",X"38",X"CD",X"0D",X"39",
		X"D8",X"FD",X"35",X"01",X"C3",X"44",X"38",X"3E",X"05",X"A2",X"20",X"F8",X"CD",X"0D",X"39",X"D8",
		X"FD",X"34",X"01",X"C3",X"D4",X"38",X"FD",X"7E",X"02",X"DD",X"BE",X"01",X"38",X"0F",X"3E",X"0A",
		X"A2",X"20",X"E1",X"CD",X"0D",X"39",X"D8",X"FD",X"35",X"02",X"C3",X"D4",X"38",X"3E",X"0A",X"A2",
		X"20",X"D2",X"CD",X"0D",X"39",X"D8",X"FD",X"34",X"02",X"C3",X"D4",X"38",X"C9",X"DD",X"21",X"96",
		X"61",X"DD",X"7E",X"00",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"27",X"5F",X"CB",
		X"27",X"83",X"06",X"00",X"4F",X"21",X"A2",X"0D",X"09",X"DD",X"7E",X"01",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"D6",X"03",X"5F",X"CB",X"3F",X"4F",X"09",X"7E",X"CB",X"43",X"28",X"0B",
		X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C3",X"4D",X"39",X"E6",X"0F",X"5F",X"A2",X"C2",
		X"54",X"39",X"37",X"C9",X"A7",X"C9",X"2A",X"99",X"61",X"23",X"22",X"99",X"61",X"7C",X"FE",X"00",
		X"28",X"13",X"FE",X"02",X"38",X"4A",X"7D",X"FE",X"58",X"38",X"45",X"21",X"00",X"00",X"22",X"99",
		X"61",X"3E",X"07",X"18",X"13",X"7D",X"FE",X"01",X"28",X"F7",X"FE",X"1E",X"20",X"04",X"3E",X"06",
		X"18",X"06",X"FE",X"B4",X"20",X"2A",X"3E",X"05",X"06",X"06",X"DD",X"21",X"9C",X"61",X"11",X"00",
		X"04",X"DD",X"6E",X"00",X"DD",X"23",X"DD",X"66",X"00",X"DD",X"23",X"4F",X"AF",X"BC",X"79",X"28",
		X"0D",X"19",X"77",X"23",X"77",X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"77",X"2B",X"77",X"10",X"E1",
		X"C9",X"21",X"AA",X"60",X"35",X"C2",X"48",X"3A",X"2A",X"63",X"60",X"3A",X"62",X"60",X"FE",X"00",
		X"28",X"04",X"36",X"06",X"18",X"02",X"36",X"05",X"3A",X"60",X"60",X"4F",X"CD",X"24",X"1D",X"22",
		X"63",X"60",X"21",X"00",X"60",X"CB",X"E6",X"21",X"61",X"60",X"34",X"7E",X"FE",X"17",X"20",X"0F",
		X"36",X"00",X"21",X"60",X"60",X"34",X"7E",X"FE",X"04",X"20",X"16",X"36",X"00",X"18",X"12",X"FE",
		X"0C",X"20",X"0E",X"3A",X"60",X"60",X"FE",X"00",X"20",X"07",X"3A",X"62",X"60",X"2F",X"32",X"62",
		X"60",X"3A",X"AB",X"60",X"32",X"AA",X"60",X"3A",X"60",X"60",X"FE",X"00",X"20",X"3A",X"3A",X"61",
		X"60",X"FE",X"01",X"28",X"1B",X"FE",X"0C",X"20",X"2F",X"06",X"04",X"11",X"05",X"00",X"21",X"2B",
		X"60",X"CB",X"46",X"20",X"05",X"19",X"10",X"F9",X"18",X"1E",X"CB",X"86",X"CB",X"CE",X"18",X"18",
		X"06",X"04",X"11",X"05",X"00",X"21",X"2B",X"60",X"CB",X"46",X"20",X"05",X"19",X"10",X"F9",X"18",
		X"07",X"E5",X"21",X"00",X"60",X"CB",X"EE",X"E1",X"21",X"CA",X"61",X"35",X"21",X"B6",X"61",X"35",
		X"23",X"20",X"22",X"2B",X"36",X"3C",X"23",X"E5",X"23",X"34",X"06",X"04",X"21",X"CE",X"61",X"AF",
		X"BE",X"28",X"01",X"35",X"23",X"10",X"F9",X"21",X"E1",X"61",X"BE",X"28",X"01",X"35",X"E1",X"7E",
		X"FE",X"F0",X"30",X"01",X"34",X"23",X"23",X"35",X"C9",X"E5",X"D5",X"F5",X"7A",X"FE",X"01",X"28",
		X"07",X"38",X"0A",X"21",X"93",X"0D",X"18",X"08",X"21",X"84",X"0D",X"18",X"03",X"21",X"7A",X"0D",
		X"F1",X"5F",X"16",X"00",X"19",X"7E",X"D1",X"E1",X"C9",X"3A",X"C9",X"61",X"E6",X"FF",X"28",X"03",
		X"C3",X"F9",X"3A",X"3A",X"26",X"60",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"98",
		X"61",X"BE",X"C0",X"FE",X"02",X"DA",X"98",X"3B",X"CA",X"61",X"3B",X"FE",X"04",X"CA",X"2E",X"3B",
		X"3A",X"27",X"60",X"D6",X"04",X"57",X"3A",X"28",X"60",X"00",X"5F",X"CD",X"0A",X"3C",X"46",X"1D",
		X"CD",X"0A",X"3C",X"7E",X"B8",X"28",X"21",X"78",X"FE",X"36",X"20",X"05",X"23",X"AF",X"C3",X"CA",
		X"3B",X"1C",X"7A",X"C6",X"08",X"57",X"CD",X"0A",X"3C",X"3E",X"35",X"BE",X"C0",X"D5",X"11",X"20",
		X"00",X"19",X"D1",X"3E",X"01",X"C3",X"CA",X"3B",X"C9",X"2A",X"CB",X"61",X"3A",X"C9",X"61",X"08",
		X"AF",X"32",X"C9",X"61",X"08",X"FE",X"02",X"28",X"0A",X"38",X"0C",X"FE",X"03",X"28",X"0C",X"3E",
		X"06",X"18",X"0A",X"3E",X"07",X"18",X"06",X"3E",X"05",X"18",X"02",X"3E",X"04",X"CD",X"EA",X"3B",
		X"CD",X"EB",X"22",X"CD",X"7B",X"46",X"21",X"5F",X"60",X"CB",X"9E",X"C3",X"A3",X"3A",X"3A",X"27",
		X"60",X"C6",X"05",X"57",X"3A",X"28",X"60",X"C6",X"05",X"5F",X"CD",X"0A",X"3C",X"7E",X"14",X"CD",
		X"0A",X"3C",X"BE",X"28",X"1B",X"3E",X"3E",X"BE",X"20",X"05",X"3E",X"03",X"C3",X"CA",X"3B",X"7B",
		X"D6",X"08",X"5F",X"CD",X"0A",X"3C",X"3E",X"3D",X"BE",X"C0",X"2B",X"3E",X"02",X"C3",X"CA",X"3B",
		X"C9",X"3A",X"27",X"60",X"C6",X"04",X"57",X"3A",X"28",X"60",X"D6",X"04",X"5F",X"CD",X"0A",X"3C",
		X"7E",X"1D",X"CD",X"0A",X"3C",X"BE",X"28",X"1F",X"3E",X"35",X"BE",X"20",X"0A",X"D5",X"11",X"20",
		X"00",X"19",X"D1",X"AF",X"C3",X"CA",X"3B",X"7A",X"D6",X"08",X"57",X"CD",X"0A",X"3C",X"3E",X"36",
		X"BE",X"C0",X"3E",X"01",X"C3",X"CA",X"3B",X"C9",X"C3",X"80",X"00",X"3C",X"57",X"3A",X"28",X"60",
		X"D6",X"03",X"5F",X"CD",X"0A",X"3C",X"7E",X"15",X"CD",X"0A",X"3C",X"BE",X"28",X"1B",X"3E",X"3D",
		X"BE",X"20",X"06",X"2B",X"3E",X"03",X"C3",X"CA",X"3B",X"7B",X"C6",X"08",X"5F",X"CD",X"0A",X"3C",
		X"3E",X"3E",X"BE",X"C0",X"3E",X"02",X"C3",X"CA",X"3B",X"C9",X"08",X"3A",X"C9",X"61",X"FE",X"00",
		X"C2",X"F9",X"3A",X"08",X"47",X"3C",X"32",X"C9",X"61",X"78",X"22",X"CB",X"61",X"08",X"3E",X"01",
		X"32",X"CA",X"61",X"08",X"CD",X"EA",X"3B",X"C3",X"FE",X"3B",X"F5",X"E5",X"06",X"01",X"7D",X"21",
		X"1D",X"0D",X"BE",X"28",X"06",X"04",X"23",X"23",X"C3",X"F2",X"3B",X"E1",X"F1",X"C9",X"CD",X"EB",
		X"22",X"CD",X"7B",X"46",X"21",X"5F",X"60",X"CB",X"9E",X"C9",X"F5",X"C5",X"7A",X"E6",X"F8",X"06",
		X"00",X"4F",X"CB",X"21",X"CB",X"10",X"CB",X"21",X"CB",X"10",X"21",X"A0",X"D0",X"09",X"7B",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"06",X"00",X"4F",X"09",X"C1",X"F1",X"C9",X"E5",X"21",X"5F",X"60",
		X"CB",X"66",X"C2",X"AE",X"3C",X"D5",X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"3A",X"9F",X"60",
		X"18",X"03",X"3A",X"A2",X"60",X"08",X"21",X"10",X"0E",X"AF",X"BB",X"20",X"15",X"08",X"06",X"00",
		X"4F",X"09",X"7E",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"06",X"00",X"0E",X"00",X"57",
		X"18",X"10",X"1D",X"CB",X"23",X"CB",X"23",X"16",X"00",X"19",X"08",X"5F",X"19",X"06",X"00",X"4E",
		X"16",X"00",X"3A",X"65",X"60",X"FE",X"00",X"20",X"06",X"DD",X"21",X"68",X"60",X"18",X"04",X"DD",
		X"21",X"6B",X"60",X"DD",X"7E",X"02",X"82",X"27",X"DD",X"77",X"02",X"DD",X"7E",X"01",X"89",X"27",
		X"DD",X"77",X"01",X"DD",X"7E",X"00",X"88",X"27",X"DD",X"77",X"00",X"3A",X"65",X"60",X"FE",X"00",
		X"20",X"05",X"21",X"C4",X"D2",X"18",X"03",X"21",X"C3",X"D2",X"CD",X"06",X"1E",X"D1",X"E1",X"C9",
		X"E5",X"D5",X"C5",X"21",X"44",X"60",X"11",X"FB",X"FF",X"06",X"06",X"AF",X"CB",X"4E",X"28",X"04",
		X"37",X"C3",X"C5",X"3C",X"A7",X"17",X"19",X"10",X"F3",X"C1",X"D1",X"E1",X"C9",X"C5",X"D5",X"E5",
		X"06",X"09",X"11",X"05",X"00",X"21",X"21",X"60",X"CB",X"86",X"CB",X"8E",X"19",X"10",X"F9",X"DD",
		X"E5",X"FD",X"E5",X"F5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"F1",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"C9",X"DD",X"21",X"43",X"0D",X"06",X"14",X"1E",X"00",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"7E",X"FE",X"36",X"20",X"03",X"A7",X"18",X"01",X"37",X"CB",X"13",X"CB",X"12",X"CB",X"11",
		X"DD",X"2B",X"DD",X"2B",X"10",X"E5",X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"21",X"A3",X"60",
		X"18",X"03",X"21",X"A6",X"60",X"73",X"23",X"72",X"23",X"71",X"C9",X"E5",X"0E",X"00",X"06",X"02",
		X"11",X"1C",X"0E",X"1A",X"13",X"BD",X"C2",X"3E",X"3D",X"1A",X"BC",X"CA",X"64",X"3D",X"13",X"10",
		X"F2",X"0C",X"06",X"0C",X"1A",X"13",X"BD",X"C2",X"4F",X"3D",X"1A",X"BC",X"CA",X"64",X"3D",X"13",
		X"10",X"F2",X"0C",X"06",X"10",X"1A",X"13",X"BD",X"C2",X"60",X"3D",X"1A",X"BC",X"CA",X"64",X"3D",
		X"13",X"10",X"F2",X"0C",X"06",X"00",X"DD",X"21",X"58",X"0E",X"CB",X"21",X"CB",X"21",X"DD",X"09",
		X"DD",X"7E",X"00",X"77",X"E5",X"11",X"00",X"04",X"19",X"36",X"02",X"E1",X"23",X"DD",X"7E",X"01",
		X"77",X"E5",X"19",X"36",X"00",X"E1",X"D5",X"11",X"E0",X"FF",X"19",X"D1",X"DD",X"7E",X"02",X"77",
		X"E5",X"19",X"36",X"00",X"E1",X"2B",X"DD",X"7E",X"03",X"77",X"19",X"36",X"00",X"E1",X"C9",X"E5",
		X"2A",X"99",X"61",X"7C",X"FE",X"00",X"20",X"09",X"7D",X"FE",X"1F",X"38",X"08",X"FE",X"B4",X"38",
		X"08",X"1E",X"01",X"18",X"06",X"1E",X"03",X"18",X"02",X"1E",X"02",X"E1",X"C9",X"D5",X"3E",X"DA",
		X"08",X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"3A",X"9F",X"60",X"18",X"03",X"3A",X"A2",X"60",
		X"FE",X"00",X"28",X"0D",X"FE",X"03",X"28",X"06",X"47",X"08",X"05",X"80",X"18",X"02",X"3E",X"DD",
		X"77",X"DD",X"21",X"26",X"60",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"00",X"8E",X"DD",X"21",X"49",
		X"60",X"DD",X"36",X"00",X"82",X"CD",X"3F",X"3E",X"3E",X"09",X"81",X"DD",X"77",X"02",X"DD",X"70",
		X"01",X"DD",X"36",X"04",X"0F",X"7B",X"FE",X"02",X"38",X"0E",X"28",X"06",X"DD",X"36",X"03",X"E0",
		X"18",X"0A",X"DD",X"36",X"03",X"DC",X"18",X"04",X"DD",X"36",X"03",X"D8",X"E5",X"21",X"00",X"60",
		X"CB",X"D6",X"06",X"1E",X"C5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"CD",X"5A",X"2D",X"C1",X"10",
		X"F3",X"AF",X"32",X"49",X"60",X"21",X"26",X"60",X"CB",X"CE",X"E1",X"36",X"FF",X"D1",X"C9",X"E5",
		X"D5",X"11",X"A0",X"D0",X"A7",X"ED",X"52",X"4D",X"3E",X"E0",X"A5",X"6F",X"06",X"02",X"CB",X"3C",
		X"CB",X"1D",X"10",X"FA",X"45",X"CB",X"21",X"CB",X"21",X"CB",X"21",X"D1",X"E1",X"C9",X"E5",X"16",
		X"00",X"FE",X"5E",X"28",X"2F",X"14",X"FE",X"5B",X"28",X"2A",X"14",X"FE",X"59",X"28",X"25",X"14",
		X"FE",X"5A",X"28",X"20",X"14",X"FE",X"5C",X"20",X"0A",X"23",X"7E",X"FE",X"66",X"38",X"15",X"14",
		X"14",X"18",X"11",X"14",X"FE",X"5D",X"28",X"0C",X"14",X"14",X"FE",X"5F",X"28",X"06",X"14",X"FE",
		X"60",X"28",X"01",X"14",X"E1",X"C9",X"FE",X"03",X"28",X"05",X"FE",X"02",X"28",X"12",X"C9",X"3A",
		X"65",X"60",X"FE",X"00",X"20",X"05",X"21",X"9D",X"60",X"18",X"16",X"21",X"A0",X"60",X"18",X"11",
		X"3A",X"65",X"60",X"FE",X"00",X"20",X"05",X"21",X"9E",X"60",X"18",X"3E",X"21",X"A1",X"60",X"18",
		X"39",X"7A",X"FE",X"00",X"20",X"04",X"CB",X"AE",X"18",X"2E",X"FE",X"01",X"20",X"04",X"CB",X"96",
		X"18",X"26",X"FE",X"02",X"20",X"04",X"CB",X"86",X"18",X"1E",X"FE",X"03",X"20",X"04",X"CB",X"8E",
		X"18",X"16",X"FE",X"04",X"20",X"04",X"CB",X"9E",X"18",X"0E",X"FE",X"05",X"20",X"04",X"CB",X"A6",
		X"18",X"06",X"FE",X"06",X"20",X"02",X"CB",X"B6",X"18",X"2F",X"7A",X"FE",X"00",X"20",X"04",X"CB",
		X"A6",X"18",X"1E",X"FE",X"01",X"20",X"04",X"CB",X"86",X"18",X"16",X"FE",X"07",X"20",X"04",X"CB",
		X"8E",X"18",X"0E",X"FE",X"08",X"20",X"04",X"CB",X"96",X"18",X"06",X"FE",X"09",X"20",X"02",X"CB",
		X"9E",X"2B",X"E5",X"CD",X"1C",X"31",X"E1",X"18",X"05",X"E5",X"CD",X"F4",X"30",X"E1",X"C9",X"CD",
		X"C7",X"1F",X"CD",X"8F",X"17",X"3A",X"03",X"60",X"FE",X"00",X"20",X"F3",X"C9",X"FD",X"21",X"9C",
		X"61",X"DD",X"21",X"91",X"60",X"CD",X"35",X"40",X"DD",X"21",X"92",X"60",X"CD",X"35",X"40",X"DD",
		X"21",X"93",X"60",X"CD",X"35",X"40",X"DD",X"21",X"94",X"60",X"CD",X"35",X"40",X"CD",X"A9",X"34",
		X"08",X"47",X"3E",X"06",X"90",X"28",X"13",X"47",X"08",X"CB",X"27",X"16",X"00",X"5F",X"21",X"A8",
		X"61",X"19",X"36",X"00",X"23",X"36",X"00",X"23",X"10",X"F8",X"C9",X"DD",X"E5",X"F5",X"D5",X"78",
		X"FE",X"0A",X"38",X"12",X"28",X"0A",X"FE",X"0B",X"20",X"2D",X"DD",X"21",X"A8",X"61",X"18",X"0A",
		X"DD",X"21",X"A2",X"61",X"18",X"04",X"DD",X"21",X"9C",X"61",X"DD",X"7E",X"01",X"FE",X"00",X"28",
		X"10",X"DD",X"23",X"DD",X"23",X"DD",X"E5",X"11",X"B4",X"61",X"7B",X"D1",X"BB",X"28",X"08",X"18",
		X"E9",X"DD",X"75",X"00",X"DD",X"74",X"01",X"D1",X"F1",X"DD",X"E1",X"C9",X"F5",X"C5",X"E5",X"AF",
		X"06",X"18",X"21",X"9C",X"61",X"77",X"23",X"10",X"FC",X"E1",X"C1",X"F1",X"C9",X"21",X"02",X"90",
		X"CB",X"6E",X"28",X"10",X"21",X"00",X"A0",X"3A",X"65",X"60",X"FE",X"00",X"20",X"04",X"CB",X"86",
		X"18",X"02",X"CB",X"C6",X"C9",X"F5",X"C5",X"D5",X"06",X"0C",X"11",X"9C",X"61",X"1A",X"BD",X"20",
		X"06",X"13",X"1A",X"1B",X"BC",X"28",X"06",X"13",X"13",X"10",X"F2",X"18",X"04",X"AF",X"12",X"13");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
