library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"12",X"D1",X"C1",X"F1",X"C9",X"06",X"06",X"DD",X"21",X"A8",X"61",X"DD",X"7E",X"01",X"FE",X"00",
		X"28",X"1C",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"E5",X"C5",X"CD",X"2B",X"3D",X"36",X"E5",
		X"21",X"A9",X"60",X"34",X"C1",X"DD",X"E1",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"23",
		X"DD",X"23",X"10",X"D7",X"C9",X"AF",X"06",X"03",X"DD",X"4E",X"00",X"CD",X"3B",X"33",X"FD",X"75",
		X"00",X"FD",X"23",X"FD",X"74",X"00",X"FD",X"23",X"3C",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"DD",
		X"23",X"10",X"E5",X"C9",X"06",X"0C",X"DD",X"21",X"9C",X"61",X"DD",X"7E",X"01",X"FE",X"00",X"28",
		X"16",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"E5",X"C5",X"CD",X"2B",X"3D",X"C1",X"DD",X"E1",
		X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"23",X"DD",X"23",X"10",X"DD",X"C9",X"3A",X"B4",
		X"61",X"E6",X"0F",X"CA",X"A4",X"40",X"21",X"21",X"60",X"CB",X"8E",X"CB",X"86",X"06",X"04",X"21",
		X"2B",X"60",X"11",X"05",X"00",X"1F",X"D2",X"9D",X"40",X"CB",X"86",X"CB",X"8E",X"19",X"10",X"F5",
		X"AF",X"32",X"B4",X"61",X"CD",X"F8",X"40",X"CD",X"B0",X"3C",X"E6",X"0F",X"28",X"1D",X"CD",X"5C",
		X"2E",X"CD",X"CC",X"40",X"06",X"04",X"21",X"2B",X"60",X"C3",X"C2",X"40",X"D5",X"11",X"05",X"00",
		X"19",X"D1",X"CB",X"4E",X"28",X"03",X"CD",X"BA",X"42",X"10",X"F1",X"C9",X"3A",X"C3",X"61",X"47",
		X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"CB",X"2F",X"5F",X"CB",X"48",X"20",X"10",X"CB",X"50",X"20",
		X"08",X"CB",X"58",X"28",X"12",X"3E",X"CC",X"18",X"06",X"3E",X"80",X"18",X"02",X"3E",X"33",X"21",
		X"B5",X"61",X"86",X"77",X"30",X"01",X"1C",X"C9",X"CD",X"26",X"1F",X"21",X"A6",X"0E",X"FE",X"33",
		X"DA",X"05",X"41",X"3E",X"32",X"5F",X"16",X"00",X"19",X"5E",X"21",X"D8",X"0E",X"3A",X"02",X"90",
		X"CB",X"4F",X"20",X"03",X"21",X"E8",X"0E",X"3A",X"B7",X"61",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"83",X"FE",X"10",X"38",X"02",X"3E",X"0F",X"5F",X"19",X"7E",X"32",X"C3",X"61",X"C9",
		X"CB",X"47",X"20",X"1B",X"CB",X"4F",X"20",X"2A",X"CB",X"57",X"20",X"39",X"3E",X"02",X"83",X"5F",
		X"CD",X"0A",X"3C",X"7E",X"FE",X"35",X"28",X"3F",X"FE",X"37",X"28",X"3B",X"C3",X"85",X"41",X"7A",
		X"D6",X"01",X"57",X"CD",X"0A",X"3C",X"7E",X"FE",X"3D",X"28",X"2C",X"FE",X"3F",X"28",X"28",X"C3",
		X"85",X"41",X"7B",X"D6",X"07",X"5F",X"CD",X"0A",X"3C",X"7E",X"FE",X"35",X"28",X"19",X"FE",X"37",
		X"28",X"15",X"C3",X"85",X"41",X"3E",X"08",X"82",X"57",X"CD",X"0A",X"3C",X"7E",X"FE",X"3F",X"28",
		X"06",X"FE",X"3D",X"28",X"02",X"A7",X"C9",X"37",X"C9",X"CB",X"47",X"20",X"2C",X"CB",X"4F",X"20",
		X"4B",X"CB",X"57",X"20",X"6A",X"3E",X"02",X"83",X"47",X"5F",X"CD",X"0A",X"3C",X"7E",X"FE",X"4A",
		X"CA",X"22",X"42",X"FE",X"45",X"28",X"7B",X"78",X"C6",X"02",X"5F",X"CD",X"0A",X"3C",X"7E",X"FE",
		X"41",X"28",X"6F",X"FE",X"46",X"28",X"6B",X"18",X"67",X"7A",X"D6",X"01",X"47",X"57",X"CD",X"0A",
		X"3C",X"7E",X"FE",X"45",X"28",X"5C",X"FE",X"46",X"28",X"58",X"78",X"D6",X"02",X"57",X"CD",X"0A",
		X"3C",X"7E",X"FE",X"4A",X"28",X"4C",X"FE",X"41",X"28",X"48",X"18",X"44",X"7B",X"D6",X"01",X"47",
		X"5F",X"CD",X"0A",X"3C",X"7E",X"FE",X"49",X"28",X"39",X"FE",X"43",X"28",X"35",X"78",X"D6",X"06",
		X"5F",X"CD",X"0A",X"3C",X"7E",X"FE",X"41",X"28",X"29",X"FE",X"46",X"28",X"25",X"18",X"21",X"3E",
		X"02",X"82",X"47",X"57",X"CD",X"0A",X"3C",X"7E",X"FE",X"44",X"28",X"16",X"FE",X"47",X"28",X"12",
		X"78",X"C6",X"06",X"57",X"CD",X"0A",X"3C",X"7E",X"FE",X"4A",X"28",X"06",X"FE",X"41",X"28",X"02",
		X"A7",X"C9",X"37",X"C9",X"DD",X"7E",X"00",X"FE",X"02",X"38",X"0A",X"28",X"0C",X"FE",X"04",X"28",
		X"0C",X"DD",X"34",X"02",X"C9",X"DD",X"35",X"01",X"C9",X"DD",X"35",X"02",X"C9",X"DD",X"34",X"01",
		X"C9",X"DD",X"21",X"BE",X"61",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"06",X"01",X"1F",X"30",X"0A",
		X"CB",X"20",X"CB",X"60",X"28",X"F7",X"AF",X"C3",X"4B",X"42",X"32",X"C8",X"61",X"C5",X"50",X"CD",
		X"11",X"39",X"C1",X"3A",X"C8",X"61",X"38",X"E8",X"32",X"C8",X"61",X"C5",X"78",X"DD",X"56",X"00",
		X"DD",X"5E",X"01",X"CD",X"30",X"41",X"C1",X"3A",X"C8",X"61",X"38",X"D4",X"50",X"C9",X"08",X"7A",
		X"E6",X"0F",X"FE",X"08",X"20",X"32",X"7B",X"E6",X"0F",X"FE",X"06",X"20",X"2B",X"08",X"E6",X"05",
		X"20",X"08",X"43",X"7A",X"CD",X"7A",X"37",X"C3",X"9F",X"42",X"42",X"7B",X"CD",X"DA",X"36",X"CB",
		X"3A",X"CB",X"1B",X"DA",X"AA",X"42",X"81",X"C3",X"9F",X"42",X"CD",X"03",X"37",X"28",X"07",X"38",
		X"07",X"CB",X"FA",X"C3",X"A6",X"42",X"37",X"C9",X"A7",X"C9",X"E5",X"D5",X"C5",X"CD",X"F0",X"43",
		X"01",X"03",X"00",X"21",X"BA",X"61",X"11",X"BD",X"61",X"ED",X"B0",X"AF",X"32",X"C1",X"61",X"32",
		X"C2",X"61",X"21",X"BD",X"61",X"7E",X"23",X"56",X"23",X"5E",X"CD",X"7E",X"42",X"D2",X"3A",X"43",
		X"CD",X"E6",X"42",X"C3",X"BA",X"43",X"DD",X"21",X"BE",X"61",X"E1",X"C1",X"C5",X"E5",X"3E",X"04",
		X"90",X"4F",X"06",X"00",X"21",X"C4",X"61",X"09",X"56",X"CD",X"11",X"39",X"38",X"13",X"D5",X"7A",
		X"21",X"BE",X"61",X"56",X"23",X"5E",X"CD",X"30",X"41",X"D1",X"38",X"05",X"21",X"BD",X"61",X"72",
		X"C9",X"3A",X"C1",X"61",X"B2",X"32",X"C1",X"61",X"21",X"BD",X"61",X"7E",X"47",X"A3",X"28",X"09",
		X"78",X"23",X"56",X"23",X"5E",X"CD",X"30",X"41",X"D0",X"3A",X"BD",X"61",X"47",X"3A",X"C1",X"61",
		X"B0",X"32",X"C1",X"61",X"CD",X"41",X"42",X"C3",X"0C",X"43",X"21",X"BD",X"61",X"7E",X"23",X"56",
		X"23",X"5E",X"CD",X"89",X"41",X"30",X"12",X"3A",X"BD",X"61",X"47",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"20",X"CB",X"20",X"B0",X"E6",X"0F",X"32",X"BD",X"61",X"21",X"BD",X"61",X"7E",X"23",X"56",X"23",
		X"5E",X"FE",X"02",X"28",X"0D",X"38",X"12",X"FE",X"04",X"28",X"0B",X"7B",X"D6",X"04",X"5F",X"C3",
		X"7B",X"43",X"1D",X"C3",X"7B",X"43",X"14",X"14",X"14",X"14",X"14",X"CD",X"0A",X"3C",X"7E",X"FE",
		X"63",X"C2",X"BA",X"43",X"CD",X"E5",X"3F",X"CD",X"2B",X"3D",X"E5",X"21",X"01",X"60",X"CB",X"FE",
		X"21",X"5F",X"60",X"CB",X"B6",X"E1",X"C1",X"C5",X"21",X"B4",X"61",X"3E",X"04",X"90",X"28",X"0B",
		X"FE",X"02",X"28",X"0C",X"38",X"0F",X"CB",X"DE",X"C3",X"CE",X"43",X"CB",X"C6",X"C3",X"CE",X"43",
		X"CB",X"D6",X"C3",X"CE",X"43",X"CB",X"CE",X"C3",X"CE",X"43",X"DD",X"21",X"BD",X"61",X"CD",X"24",
		X"42",X"21",X"C2",X"61",X"34",X"7E",X"C1",X"D1",X"D5",X"C5",X"BB",X"C2",X"D2",X"42",X"C1",X"D1",
		X"E1",X"E5",X"D5",X"C5",X"3A",X"BD",X"61",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",
		X"CF",X"77",X"3A",X"BE",X"61",X"23",X"77",X"3A",X"BF",X"61",X"23",X"77",X"C1",X"D1",X"E1",X"C9",
		X"11",X"BA",X"61",X"7E",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"12",X"13",X"23",X"7E",
		X"12",X"13",X"23",X"7E",X"12",X"C9",X"11",X"05",X"00",X"06",X"04",X"21",X"2B",X"60",X"E5",X"C5",
		X"CB",X"46",X"C2",X"7A",X"44",X"19",X"10",X"F8",X"C1",X"E1",X"CB",X"4E",X"28",X"23",X"19",X"10",
		X"F9",X"21",X"5F",X"60",X"CB",X"76",X"C0",X"DD",X"21",X"21",X"60",X"DD",X"36",X"00",X"82",X"DD",
		X"36",X"01",X"58",X"DD",X"36",X"02",X"86",X"CD",X"7F",X"1F",X"DD",X"77",X"03",X"DD",X"70",X"04",
		X"C9",X"E5",X"C5",X"06",X"04",X"21",X"2B",X"60",X"CB",X"4E",X"28",X"1B",X"E5",X"DD",X"E1",X"3E",
		X"58",X"DD",X"BE",X"01",X"20",X"11",X"3E",X"86",X"DD",X"BE",X"02",X"38",X"0A",X"3E",X"94",X"DD",
		X"BE",X"02",X"30",X"03",X"C1",X"E1",X"C9",X"19",X"10",X"DE",X"C1",X"78",X"D6",X"04",X"ED",X"44",
		X"4F",X"CD",X"61",X"30",X"E1",X"CB",X"8E",X"CB",X"C6",X"C9",X"C1",X"E1",X"C9",X"3A",X"5F",X"60",
		X"CB",X"5F",X"CA",X"9A",X"44",X"ED",X"4B",X"D3",X"61",X"ED",X"5B",X"D5",X"61",X"26",X"62",X"3A",
		X"D7",X"61",X"FE",X"00",X"CA",X"CA",X"44",X"C3",X"42",X"45",X"CD",X"C4",X"45",X"01",X"CF",X"62",
		X"11",X"FF",X"62",X"3E",X"FF",X"02",X"12",X"21",X"26",X"60",X"CB",X"4E",X"C8",X"23",X"D5",X"C5",
		X"56",X"23",X"5E",X"3E",X"35",X"BB",X"DA",X"BC",X"44",X"C1",X"D1",X"C9",X"CD",X"DC",X"45",X"C1",
		X"D1",X"0D",X"02",X"26",X"62",X"6F",X"7E",X"F6",X"0F",X"77",X"0A",X"FE",X"FF",X"CA",X"3C",X"45",
		X"6F",X"CB",X"7E",X"28",X"12",X"E5",X"D5",X"11",X"F0",X"FF",X"19",X"D1",X"7E",X"E6",X"0F",X"20",
		X"05",X"CB",X"CE",X"1D",X"7D",X"12",X"E1",X"CB",X"76",X"28",X"0D",X"E5",X"2C",X"7E",X"E6",X"0F",
		X"20",X"05",X"CB",X"C6",X"1D",X"7D",X"12",X"E1",X"CB",X"6E",X"28",X"12",X"E5",X"D5",X"11",X"10",
		X"00",X"19",X"D1",X"7E",X"E6",X"0F",X"20",X"05",X"CB",X"DE",X"1D",X"7D",X"12",X"E1",X"CB",X"66",
		X"28",X"0D",X"E5",X"2D",X"7E",X"E6",X"0F",X"20",X"05",X"CB",X"D6",X"1D",X"7D",X"12",X"E1",X"0C",
		X"E5",X"21",X"01",X"90",X"CB",X"7E",X"E1",X"CA",X"CA",X"44",X"21",X"5F",X"60",X"CB",X"DE",X"ED",
		X"43",X"D3",X"61",X"ED",X"53",X"D5",X"61",X"AF",X"32",X"D7",X"61",X"C9",X"1A",X"FE",X"FF",X"CA",
		X"BE",X"45",X"1A",X"FE",X"FF",X"CA",X"B8",X"45",X"6F",X"CB",X"7E",X"28",X"12",X"E5",X"D5",X"11",
		X"F0",X"FF",X"19",X"D1",X"7E",X"E6",X"0F",X"20",X"05",X"CB",X"CE",X"0D",X"7D",X"02",X"E1",X"CB",
		X"76",X"28",X"0D",X"E5",X"2C",X"7E",X"E6",X"0F",X"20",X"05",X"CB",X"C6",X"0D",X"7D",X"02",X"E1",
		X"CB",X"6E",X"28",X"12",X"E5",X"D5",X"11",X"10",X"00",X"19",X"D1",X"7E",X"E6",X"0F",X"20",X"05",
		X"CB",X"DE",X"0D",X"7D",X"02",X"E1",X"CB",X"66",X"28",X"0D",X"E5",X"2D",X"7E",X"E6",X"0F",X"20",
		X"05",X"CB",X"D6",X"0D",X"7D",X"02",X"E1",X"1C",X"E5",X"21",X"01",X"90",X"CB",X"7E",X"E1",X"CA",
		X"42",X"45",X"21",X"5F",X"60",X"CB",X"DE",X"ED",X"43",X"D3",X"61",X"ED",X"53",X"D5",X"61",X"CB",
		X"C7",X"32",X"D7",X"61",X"C9",X"C3",X"42",X"45",X"0A",X"FE",X"FF",X"C2",X"CA",X"44",X"21",X"5F",
		X"60",X"CB",X"9E",X"C9",X"11",X"10",X"00",X"21",X"00",X"62",X"E5",X"06",X"0B",X"7E",X"E6",X"F0",
		X"77",X"23",X"10",X"F9",X"E1",X"19",X"3E",X"B0",X"BD",X"20",X"EF",X"C9",X"CB",X"3A",X"CB",X"3A",
		X"CB",X"3A",X"CB",X"3A",X"7B",X"D6",X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"4F",
		X"3E",X"0A",X"91",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"B2",X"C9",X"DD",X"21",X"A2",
		X"0D",X"21",X"A0",X"62",X"06",X"0B",X"11",X"F0",X"FF",X"E5",X"C5",X"06",X"05",X"DD",X"7E",X"00",
		X"4F",X"E6",X"0F",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"77",X"19",X"79",X"E6",X"F0",
		X"77",X"19",X"DD",X"23",X"10",X"E7",X"DD",X"7E",X"00",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"77",X"C1",X"E1",X"DD",X"23",X"23",X"10",X"D0",X"C9",X"11",X"C4",X"46",X"DD",X"21",X"1D",
		X"0D",X"3E",X"01",X"01",X"F0",X"FF",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"F5",X"7E",X"FE",X"36",
		X"21",X"00",X"62",X"1A",X"6F",X"28",X"0D",X"CB",X"A6",X"2B",X"CB",X"B6",X"09",X"CB",X"B6",X"23",
		X"CB",X"A6",X"18",X"0B",X"CB",X"BE",X"2B",X"CB",X"BE",X"09",X"CB",X"AE",X"23",X"CB",X"AE",X"F1",
		X"13",X"DD",X"23",X"DD",X"23",X"3C",X"FE",X"15",X"20",X"CC",X"C9",X"E5",X"21",X"C4",X"46",X"05",
		X"48",X"06",X"00",X"09",X"EB",X"01",X"F0",X"FF",X"E1",X"7E",X"32",X"C8",X"61",X"FE",X"36",X"21",
		X"00",X"62",X"1A",X"6F",X"28",X"1A",X"3A",X"C8",X"61",X"FE",X"3E",X"C0",X"CB",X"FE",X"CB",X"A6",
		X"2B",X"CB",X"FE",X"CB",X"B6",X"09",X"CB",X"EE",X"CB",X"B6",X"23",X"CB",X"EE",X"CB",X"A6",X"C9",
		X"CB",X"E6",X"CB",X"BE",X"2B",X"CB",X"F6",X"CB",X"BE",X"09",X"CB",X"F6",X"CB",X"AE",X"23",X"CB",
		X"E6",X"CB",X"AE",X"C9",X"31",X"A2",X"72",X"12",X"63",X"33",X"94",X"74",X"44",X"24",X"97",X"77",
		X"47",X"27",X"68",X"38",X"A9",X"79",X"19",X"3A",X"CD",X"26",X"1F",X"FE",X"1E",X"38",X"02",X"3E",
		X"1E",X"21",X"88",X"47",X"32",X"C8",X"61",X"3D",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"21",
		X"A6",X"47",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"47",X"F5",X"3A",X"B8",X"61",X"4F",X"78",
		X"06",X"00",X"17",X"38",X"03",X"04",X"18",X"FA",X"C5",X"79",X"07",X"10",X"FD",X"C1",X"CB",X"3F",
		X"10",X"FC",X"47",X"F1",X"B8",X"20",X"3C",X"3A",X"B6",X"61",X"FE",X"3B",X"20",X"35",X"21",X"D2",
		X"61",X"7E",X"34",X"E6",X"03",X"21",X"CE",X"61",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"FE",
		X"00",X"20",X"20",X"E5",X"21",X"AE",X"47",X"3A",X"02",X"90",X"CB",X"47",X"20",X"03",X"21",X"CD",
		X"47",X"3A",X"B7",X"61",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"85",X"6F",X"3E",X"00",X"8C",X"67",
		X"7E",X"E1",X"77",X"FD",X"21",X"C4",X"61",X"11",X"05",X"00",X"DD",X"21",X"2C",X"60",X"21",X"CE",
		X"61",X"06",X"04",X"7E",X"FE",X"00",X"28",X"18",X"D5",X"DD",X"56",X"00",X"DD",X"5E",X"01",X"CD",
		X"DC",X"45",X"5F",X"16",X"62",X"1A",X"E6",X"0F",X"D1",X"FE",X"0F",X"28",X"03",X"FD",X"77",X"00",
		X"FD",X"23",X"DD",X"19",X"23",X"10",X"DC",X"C9",X"00",X"02",X"03",X"04",X"01",X"02",X"03",X"02",
		X"03",X"04",X"03",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"05",X"05",X"05",X"04",X"03",X"02",X"01",X"01",X"03",X"03",
		X"04",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"08",X"08",X"09",X"09",X"0A",X"0A",X"0B",X"0B",
		X"0C",X"0C",X"0D",X"0D",X"0E",X"0E",X"0F",X"0F",X"10",X"10",X"11",X"11",X"12",X"0A",X"0B",X"0C",
		X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"1A",X"1B",X"1C",
		X"1D",X"1E",X"1F",X"20",X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"F5",X"E5",X"D5",X"C5",
		X"DD",X"E5",X"06",X"0C",X"21",X"9D",X"D0",X"11",X"20",X"00",X"3E",X"FF",X"77",X"23",X"77",X"19",
		X"77",X"2B",X"77",X"19",X"10",X"F6",X"06",X"0C",X"21",X"9D",X"D4",X"3E",X"01",X"77",X"23",X"77",
		X"19",X"77",X"2B",X"77",X"19",X"10",X"F6",X"06",X"16",X"21",X"9E",X"D0",X"DD",X"21",X"08",X"49",
		X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",X"F7",X"06",X"13",X"21",X"9D",X"D0",X"DD",X"21",
		X"1E",X"49",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",X"10",X"F7",X"DD",X"E1",X"C1",X"D1",X"E1",
		X"F1",X"C9",X"CD",X"EC",X"47",X"E5",X"D5",X"C5",X"F5",X"E5",X"D5",X"C5",X"F5",X"11",X"DE",X"D0",
		X"06",X"05",X"21",X"01",X"00",X"39",X"3E",X"00",X"ED",X"6F",X"CD",X"B2",X"48",X"ED",X"6F",X"CD",
		X"C0",X"48",X"23",X"10",X"F1",X"F1",X"C1",X"D1",X"E1",X"F1",X"C1",X"D1",X"E1",X"C5",X"D5",X"E5",
		X"DD",X"E5",X"FD",X"E5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"11",X"5D",X"D3",X"06",X"03",
		X"21",X"00",X"00",X"39",X"3E",X"00",X"ED",X"67",X"CD",X"CE",X"48",X"ED",X"67",X"CD",X"CE",X"48",
		X"23",X"ED",X"67",X"CD",X"CE",X"48",X"ED",X"67",X"CD",X"DE",X"48",X"23",X"10",X"E6",X"FD",X"E1",
		X"DD",X"E1",X"E1",X"D1",X"C1",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"C9",X"76",X"CD",X"D5",
		X"22",X"C9",X"E5",X"F5",X"6B",X"62",X"77",X"11",X"20",X"00",X"19",X"5D",X"54",X"F1",X"E1",X"C9",
		X"E5",X"F5",X"6B",X"62",X"77",X"11",X"80",X"00",X"19",X"5D",X"54",X"F1",X"E1",X"C9",X"E5",X"F5",
		X"6B",X"62",X"77",X"11",X"20",X"00",X"A7",X"ED",X"52",X"5D",X"54",X"F1",X"E1",X"C9",X"E5",X"F5",
		X"6B",X"62",X"77",X"11",X"A0",X"00",X"A7",X"ED",X"52",X"5D",X"54",X"F1",X"E1",X"C9",X"21",X"00",
		X"60",X"7E",X"CD",X"42",X"48",X"DD",X"21",X"00",X"90",X"DD",X"CB",X"00",X"76",X"20",X"FA",X"DD",
		X"CB",X"00",X"76",X"28",X"FA",X"23",X"18",X"E9",X"0A",X"2A",X"FF",X"FF",X"FF",X"0C",X"2A",X"FF",
		X"FF",X"FF",X"0B",X"2A",X"FF",X"FF",X"FF",X"0E",X"2A",X"FF",X"FF",X"FF",X"0D",X"2A",X"11",X"15",
		X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"12",X"21",X"2A",X"FF",X"FF",X"FF",X"FF",X"FF",X"12",X"22",
		X"2A",X"36",X"0D",X"19",X"36",X"FF",X"19",X"C3",X"EB",X"1D",X"36",X"1D",X"19",X"36",X"FF",X"19",
		X"C3",X"FE",X"1D",X"D5",X"AF",X"32",X"E0",X"61",X"C3",X"6E",X"37",X"3A",X"26",X"60",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"C3",X"77",X"36",X"32",X"5F",X"60",X"32",X"E3",X"61",X"C3",X"DC",X"02",
		X"21",X"5E",X"60",X"35",X"35",X"21",X"E2",X"61",X"34",X"C3",X"E1",X"03",X"32",X"65",X"60",X"21",
		X"E3",X"61",X"7E",X"FE",X"00",X"CA",X"86",X"49",X"3A",X"5F",X"60",X"CB",X"4F",X"CA",X"81",X"49",
		X"35",X"35",X"AF",X"32",X"E2",X"61",X"C3",X"E5",X"03",X"21",X"E3",X"61",X"34",X"CD",X"2F",X"3F",
		X"C3",X"45",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"19",X"58",X"A0",X"00",X"41",X"19",X"60",X"1C",X"06",X"21",X"11",X"68",X"A4",X"F6",X"5A",
		X"01",X"44",X"04",X"80",X"09",X"A1",X"00",X"A0",X"05",X"01",X"00",X"00",X"40",X"22",X"00",X"00",
		X"02",X"10",X"A0",X"00",X"04",X"00",X"00",X"29",X"01",X"20",X"01",X"04",X"85",X"0D",X"21",X"33",
		X"9B",X"1F",X"02",X"1E",X"C9",X"C0",X"88",X"84",X"84",X"4A",X"80",X"C2",X"42",X"14",X"C6",X"46",
		X"46",X"00",X"D0",X"A4",X"A1",X"4C",X"C2",X"99",X"18",X"8A",X"42",X"E8",X"42",X"13",X"C8",X"E0",
		X"11",X"10",X"18",X"62",X"22",X"40",X"41",X"02",X"80",X"04",X"50",X"08",X"18",X"10",X"40",X"80",
		X"F0",X"20",X"A0",X"00",X"0D",X"04",X"00",X"00",X"14",X"60",X"80",X"40",X"00",X"10",X"04",X"60",
		X"10",X"16",X"58",X"87",X"71",X"15",X"01",X"92",X"A5",X"01",X"06",X"02",X"02",X"01",X"00",X"C0",
		X"23",X"01",X"10",X"85",X"81",X"80",X"50",X"22",X"44",X"0B",X"19",X"02",X"8B",X"B5",X"AF",X"AC",
		X"00",X"00",X"00",X"82",X"80",X"24",X"00",X"10",X"00",X"00",X"01",X"50",X"00",X"80",X"10",X"80",
		X"20",X"00",X"09",X"04",X"01",X"00",X"40",X"00",X"00",X"00",X"12",X"00",X"A0",X"81",X"22",X"63",
		X"5B",X"4E",X"0D",X"58",X"44",X"C2",X"93",X"11",X"94",X"C4",X"82",X"41",X"40",X"00",X"40",X"FA",
		X"66",X"8B",X"50",X"C5",X"2B",X"81",X"0F",X"07",X"42",X"85",X"80",X"06",X"1A",X"48",X"47",X"89",
		X"08",X"0C",X"00",X"C8",X"00",X"10",X"44",X"00",X"10",X"00",X"00",X"00",X"08",X"00",X"08",X"44",
		X"92",X"00",X"10",X"40",X"80",X"01",X"10",X"0A",X"00",X"02",X"42",X"00",X"AA",X"00",X"10",X"60",
		X"B1",X"90",X"14",X"68",X"A3",X"80",X"85",X"12",X"96",X"0A",X"02",X"10",X"21",X"05",X"81",X"03",
		X"20",X"70",X"00",X"00",X"44",X"11",X"09",X"0D",X"61",X"01",X"9A",X"A8",X"45",X"B8",X"9C",X"A7",
		X"A0",X"C2",X"83",X"21",X"40",X"20",X"20",X"00",X"08",X"20",X"81",X"00",X"35",X"08",X"00",X"90",
		X"B0",X"00",X"00",X"00",X"00",X"28",X"41",X"00",X"20",X"20",X"04",X"10",X"AC",X"84",X"A6",X"38",
		X"42",X"62",X"A2",X"2C",X"95",X"84",X"91",X"C3",X"C0",X"04",X"42",X"01",X"59",X"44",X"83",X"C0",
		X"4A",X"64",X"64",X"30",X"C0",X"2E",X"58",X"C8",X"B9",X"C3",X"E8",X"E1",X"84",X"5A",X"05",X"CE",
		X"00",X"80",X"00",X"10",X"00",X"00",X"08",X"40",X"72",X"04",X"40",X"08",X"40",X"00",X"00",X"90",
		X"01",X"00",X"00",X"00",X"01",X"40",X"00",X"00",X"90",X"A0",X"00",X"A2",X"00",X"80",X"90",X"00",
		X"74",X"80",X"29",X"01",X"F0",X"30",X"B1",X"A1",X"21",X"31",X"35",X"1D",X"09",X"1D",X"A5",X"07",
		X"21",X"F0",X"22",X"20",X"27",X"A1",X"01",X"82",X"C0",X"08",X"A4",X"11",X"38",X"B5",X"C8",X"A5",
		X"22",X"00",X"00",X"03",X"30",X"E1",X"A0",X"01",X"00",X"00",X"08",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"41",X"80",X"40",X"80",X"01",X"00",X"08",X"50",X"82",X"20",X"9F",X"4D",
		X"72",X"A9",X"06",X"4E",X"38",X"40",X"80",X"2E",X"04",X"A6",X"83",X"30",X"24",X"02",X"08",X"00",
		X"40",X"30",X"C2",X"20",X"62",X"64",X"E8",X"62",X"E8",X"DA",X"03",X"9B",X"08",X"51",X"46",X"16",
		X"88",X"14",X"00",X"22",X"05",X"C0",X"00",X"00",X"11",X"00",X"02",X"00",X"80",X"A0",X"40",X"00",
		X"00",X"01",X"00",X"02",X"00",X"08",X"80",X"11",X"00",X"00",X"1E",X"02",X"A0",X"22",X"10",X"00",
		X"43",X"E0",X"41",X"71",X"40",X"05",X"14",X"80",X"9C",X"20",X"AF",X"3B",X"4A",X"F8",X"01",X"33",
		X"31",X"02",X"51",X"A0",X"18",X"7C",X"80",X"33",X"25",X"00",X"1C",X"24",X"3E",X"EC",X"78",X"5F",
		X"21",X"00",X"00",X"11",X"04",X"04",X"01",X"00",X"00",X"04",X"00",X"00",X"10",X"00",X"00",X"14",
		X"80",X"20",X"40",X"20",X"20",X"16",X"00",X"90",X"08",X"04",X"00",X"10",X"23",X"40",X"08",X"09",
		X"C8",X"8A",X"C8",X"C8",X"CA",X"82",X"82",X"52",X"4A",X"C0",X"0A",X"4A",X"8A",X"C0",X"02",X"4A",
		X"4A",X"CA",X"C0",X"CA",X"C8",X"CA",X"CA",X"88",X"48",X"4A",X"4A",X"4A",X"4A",X"62",X"02",X"C0",
		X"DA",X"CA",X"08",X"EA",X"CA",X"4A",X"CA",X"EA",X"CA",X"8A",X"CA",X"C0",X"08",X"CA",X"82",X"88",
		X"80",X"C8",X"CA",X"C8",X"42",X"8A",X"C2",X"8A",X"8A",X"08",X"CA",X"CA",X"40",X"CA",X"C8",X"9A",
		X"30",X"34",X"15",X"34",X"25",X"35",X"24",X"25",X"10",X"10",X"35",X"15",X"20",X"35",X"31",X"15",
		X"10",X"35",X"35",X"34",X"74",X"34",X"11",X"14",X"20",X"34",X"04",X"31",X"34",X"35",X"35",X"25",
		X"2D",X"25",X"15",X"14",X"34",X"34",X"35",X"01",X"35",X"05",X"35",X"24",X"35",X"35",X"35",X"35",
		X"33",X"35",X"15",X"31",X"15",X"35",X"35",X"15",X"31",X"35",X"34",X"35",X"34",X"15",X"3D",X"35",
		X"CA",X"C0",X"CA",X"CA",X"88",X"88",X"CA",X"8A",X"4A",X"C8",X"C8",X"C2",X"C2",X"C8",X"4A",X"4A",
		X"00",X"CA",X"4A",X"CA",X"80",X"4A",X"CA",X"CA",X"42",X"C8",X"CA",X"42",X"4A",X"0A",X"40",X"CA",
		X"CA",X"CA",X"5A",X"CA",X"CA",X"CA",X"CA",X"4A",X"8A",X"A8",X"02",X"4A",X"CA",X"8A",X"4A",X"42",
		X"C2",X"8A",X"0A",X"C2",X"CA",X"4A",X"CA",X"CA",X"48",X"C2",X"88",X"CA",X"CA",X"C8",X"C2",X"C2",
		X"04",X"14",X"31",X"35",X"30",X"34",X"20",X"35",X"31",X"34",X"34",X"34",X"34",X"31",X"11",X"34",
		X"25",X"31",X"35",X"35",X"30",X"30",X"10",X"14",X"34",X"31",X"04",X"30",X"34",X"35",X"15",X"21",
		X"31",X"15",X"30",X"00",X"34",X"35",X"31",X"30",X"04",X"11",X"04",X"34",X"14",X"24",X"15",X"35",
		X"25",X"24",X"15",X"01",X"35",X"15",X"35",X"35",X"35",X"05",X"35",X"35",X"35",X"35",X"25",X"31",
		X"DA",X"88",X"40",X"9A",X"C2",X"CA",X"48",X"CA",X"CA",X"48",X"42",X"C0",X"0A",X"48",X"CA",X"C0",
		X"08",X"C2",X"42",X"CA",X"C8",X"42",X"C0",X"4A",X"C2",X"4A",X"48",X"CA",X"4A",X"E8",X"42",X"CA",
		X"C2",X"CA",X"CA",X"C2",X"8E",X"8A",X"C8",X"8A",X"4A",X"CA",X"CA",X"8A",X"8A",X"CA",X"CA",X"4A",
		X"C8",X"CA",X"C2",X"80",X"C8",X"4A",X"5A",X"42",X"C2",X"C0",X"8A",X"0A",X"80",X"CA",X"CA",X"C2",
		X"35",X"31",X"31",X"31",X"25",X"00",X"11",X"35",X"15",X"11",X"15",X"31",X"31",X"11",X"04",X"25",
		X"05",X"15",X"35",X"71",X"25",X"25",X"30",X"31",X"34",X"15",X"11",X"15",X"25",X"35",X"35",X"11",
		X"3C",X"25",X"35",X"35",X"35",X"35",X"55",X"15",X"25",X"31",X"31",X"14",X"35",X"3C",X"24",X"35",
		X"34",X"25",X"35",X"25",X"31",X"25",X"35",X"31",X"25",X"35",X"35",X"14",X"3D",X"25",X"35",X"B5",
		X"C8",X"CA",X"8A",X"CA",X"4A",X"CA",X"00",X"C8",X"0A",X"00",X"8A",X"CA",X"E2",X"82",X"CA",X"C0",
		X"CA",X"C2",X"48",X"CA",X"0A",X"CA",X"CA",X"C8",X"C8",X"88",X"8A",X"C8",X"C2",X"4A",X"42",X"0A",
		X"CA",X"CA",X"9A",X"CA",X"88",X"C2",X"CA",X"C2",X"CA",X"8A",X"CA",X"C2",X"82",X"CA",X"4A",X"CA",
		X"CA",X"C2",X"DA",X"44",X"CA",X"C8",X"CE",X"0A",X"C8",X"CA",X"48",X"0A",X"02",X"EA",X"C8",X"48",
		X"35",X"01",X"34",X"15",X"01",X"35",X"05",X"31",X"15",X"25",X"15",X"35",X"35",X"15",X"01",X"05",
		X"35",X"34",X"35",X"35",X"15",X"34",X"35",X"21",X"21",X"30",X"31",X"31",X"35",X"A5",X"15",X"31",
		X"30",X"34",X"01",X"B5",X"35",X"21",X"35",X"34",X"13",X"35",X"31",X"15",X"35",X"21",X"35",X"35",
		X"15",X"00",X"35",X"35",X"25",X"35",X"54",X"31",X"25",X"35",X"35",X"30",X"39",X"1D",X"35",X"15",
		X"88",X"80",X"C8",X"4A",X"80",X"CA",X"48",X"82",X"CA",X"C8",X"CA",X"C2",X"42",X"CA",X"C8",X"8A",
		X"88",X"42",X"8A",X"8A",X"C0",X"40",X"C2",X"CA",X"42",X"CA",X"CA",X"C2",X"0A",X"88",X"4A",X"4A",
		X"82",X"CA",X"C6",X"CA",X"08",X"8A",X"8A",X"C2",X"CA",X"CA",X"C8",X"CA",X"C2",X"CA",X"4A",X"CA",
		X"CA",X"C8",X"CA",X"8A",X"CA",X"CA",X"DA",X"C8",X"CA",X"88",X"02",X"CA",X"8A",X"4A",X"CA",X"80",
		X"10",X"24",X"14",X"24",X"15",X"11",X"25",X"11",X"01",X"01",X"34",X"30",X"3D",X"05",X"14",X"31",
		X"34",X"25",X"04",X"24",X"34",X"35",X"14",X"35",X"74",X"35",X"31",X"34",X"34",X"35",X"35",X"31",
		X"35",X"10",X"05",X"15",X"95",X"15",X"14",X"14",X"35",X"35",X"35",X"00",X"35",X"17",X"30",X"3D",
		X"05",X"24",X"05",X"35",X"25",X"25",X"24",X"3D",X"35",X"71",X"34",X"01",X"14",X"35",X"35",X"3C",
		X"8A",X"C2",X"CA",X"CA",X"C0",X"C8",X"40",X"C8",X"CA",X"C2",X"4A",X"C2",X"C2",X"CA",X"80",X"00",
		X"CA",X"C6",X"08",X"CA",X"4A",X"C8",X"80",X"C8",X"C2",X"CA",X"CA",X"88",X"C2",X"C8",X"CA",X"CA",
		X"CA",X"CA",X"CA",X"CA",X"C2",X"CA",X"C8",X"CA",X"CA",X"CA",X"CA",X"C2",X"CA",X"CA",X"CA",X"CA",
		X"C2",X"CA",X"CA",X"C2",X"DA",X"4A",X"CA",X"CA",X"CA",X"8A",X"C2",X"C0",X"CA",X"6A",X"CA",X"C2",
		X"24",X"15",X"11",X"34",X"35",X"35",X"35",X"05",X"25",X"11",X"01",X"21",X"25",X"21",X"15",X"21",
		X"25",X"11",X"11",X"35",X"15",X"35",X"34",X"31",X"35",X"31",X"14",X"34",X"35",X"35",X"35",X"35",
		X"34",X"11",X"35",X"35",X"15",X"15",X"14",X"21",X"25",X"35",X"31",X"34",X"34",X"31",X"34",X"3D",
		X"35",X"31",X"11",X"31",X"34",X"31",X"34",X"05",X"35",X"15",X"21",X"11",X"35",X"BD",X"B5",X"B4",
		X"C8",X"88",X"CA",X"8A",X"88",X"C8",X"CA",X"4A",X"4A",X"C8",X"CA",X"02",X"CA",X"C8",X"CA",X"C8",
		X"CA",X"CA",X"CA",X"40",X"C2",X"CA",X"4A",X"8A",X"CA",X"CA",X"48",X"8A",X"0A",X"CA",X"4A",X"E0",
		X"CA",X"C2",X"4A",X"CA",X"CA",X"CA",X"8A",X"C2",X"CA",X"CA",X"CA",X"08",X"8A",X"DA",X"82",X"4A",
		X"0A",X"C2",X"02",X"48",X"CA",X"CA",X"CA",X"0A",X"0A",X"C2",X"C2",X"88",X"C2",X"42",X"CA",X"42",
		X"14",X"30",X"14",X"34",X"31",X"21",X"31",X"25",X"27",X"14",X"35",X"31",X"24",X"24",X"35",X"31",
		X"04",X"25",X"B4",X"15",X"25",X"31",X"30",X"34",X"21",X"25",X"24",X"00",X"35",X"35",X"35",X"A5",
		X"B5",X"14",X"01",X"31",X"34",X"35",X"24",X"21",X"35",X"34",X"25",X"31",X"35",X"11",X"14",X"35",
		X"35",X"34",X"30",X"35",X"24",X"05",X"30",X"35",X"35",X"05",X"35",X"21",X"15",X"35",X"15",X"35",
		X"C0",X"CA",X"C2",X"C2",X"CA",X"C8",X"0A",X"C8",X"4A",X"40",X"02",X"42",X"C2",X"C8",X"CA",X"C2",
		X"4A",X"CA",X"C8",X"8A",X"42",X"8A",X"C8",X"4A",X"08",X"CA",X"C2",X"40",X"48",X"C8",X"0A",X"CA",
		X"CA",X"8A",X"4A",X"C2",X"CA",X"C2",X"CA",X"CA",X"4A",X"CA",X"C2",X"8A",X"42",X"C2",X"C2",X"C8",
		X"8E",X"8A",X"8A",X"CA",X"8A",X"C8",X"8A",X"EA",X"8A",X"02",X"02",X"C2",X"C2",X"4A",X"0A",X"C8",
		X"31",X"25",X"14",X"21",X"14",X"01",X"34",X"35",X"05",X"35",X"11",X"04",X"25",X"15",X"34",X"25",
		X"30",X"35",X"75",X"25",X"35",X"05",X"35",X"21",X"11",X"01",X"04",X"34",X"14",X"35",X"34",X"35",
		X"35",X"15",X"35",X"31",X"34",X"11",X"34",X"14",X"35",X"35",X"35",X"25",X"35",X"31",X"34",X"15",
		X"35",X"15",X"25",X"25",X"11",X"35",X"31",X"25",X"15",X"15",X"35",X"25",X"31",X"35",X"3D",X"3D",
		X"C3",X"60",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"C1",X"54",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"1B",X"56",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"AF",X"57",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"BF",X"58",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"A6",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"F1",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"FB",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"30",X"68",X"06",X"10",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"68",X"CB",X"1A",
		X"11",X"68",X"60",X"3A",X"65",X"60",X"A7",X"28",X"03",X"11",X"6B",X"60",X"CD",X"A4",X"50",X"D4",
		X"F6",X"50",X"3A",X"5F",X"60",X"C3",X"C0",X"5E",X"11",X"6B",X"60",X"3A",X"65",X"60",X"A7",X"28",
		X"03",X"11",X"68",X"60",X"C3",X"D0",X"5E",X"D8",X"3A",X"65",X"60",X"A7",X"28",X"02",X"3E",X"FF",
		X"2F",X"32",X"65",X"60",X"47",X"3A",X"02",X"90",X"E6",X"20",X"28",X"04",X"78",X"32",X"00",X"A0",
		X"C3",X"E0",X"5E",X"C9",X"21",X"73",X"60",X"01",X"00",X"09",X"C5",X"D5",X"E5",X"CD",X"2C",X"5D",
		X"30",X"0C",X"E1",X"01",X"03",X"00",X"09",X"D1",X"C1",X"0C",X"10",X"EE",X"37",X"C9",X"E1",X"D1",
		X"C1",X"DD",X"21",X"00",X"68",X"DD",X"36",X"00",X"5C",X"DD",X"36",X"01",X"4E",X"DD",X"36",X"02",
		X"0A",X"3A",X"02",X"90",X"E6",X"04",X"20",X"04",X"DD",X"36",X"02",X"03",X"DD",X"36",X"03",X"00",
		X"DD",X"71",X"04",X"EB",X"11",X"05",X"68",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"06",X"0A",X"36",
		X"FF",X"23",X"10",X"FB",X"A7",X"C9",X"FD",X"21",X"12",X"68",X"FD",X"36",X"00",X"82",X"FD",X"36",
		X"01",X"58",X"FD",X"36",X"02",X"36",X"21",X"85",X"D0",X"01",X"18",X"1A",X"CD",X"52",X"5D",X"21",
		X"4E",X"54",X"CD",X"36",X"5D",X"21",X"59",X"54",X"CD",X"36",X"5D",X"21",X"65",X"54",X"CD",X"36",
		X"5D",X"DD",X"7E",X"04",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"6F",X"54",X"19",X"EB",X"D5",
		X"21",X"DE",X"D1",X"01",X"06",X"03",X"CD",X"3F",X"5D",X"D1",X"21",X"DD",X"D0",X"01",X"07",X"03",
		X"CD",X"3F",X"5D",X"CD",X"6D",X"5D",X"CD",X"BC",X"5D",X"01",X"0A",X"05",X"21",X"E7",X"D0",X"11",
		X"20",X"00",X"C5",X"E5",X"36",X"31",X"19",X"36",X"31",X"19",X"36",X"33",X"19",X"19",X"10",X"F4",
		X"E1",X"23",X"23",X"C1",X"0D",X"20",X"EB",X"3E",X"0A",X"06",X"03",X"21",X"98",X"D1",X"CD",X"15",
		X"54",X"01",X"04",X"05",X"21",X"16",X"D1",X"C5",X"E5",X"CD",X"15",X"54",X"E1",X"2B",X"2B",X"C1",
		X"0D",X"20",X"F4",X"06",X"03",X"CD",X"15",X"54",X"3E",X"01",X"06",X"02",X"CD",X"15",X"54",X"06",
		X"05",X"21",X"0C",X"D1",X"CD",X"15",X"54",X"06",X"02",X"21",X"0A",X"D1",X"CD",X"15",X"54",X"3E",
		X"27",X"06",X"01",X"CD",X"15",X"54",X"3E",X"28",X"06",X"01",X"CD",X"15",X"54",X"3E",X"24",X"06",
		X"01",X"CD",X"15",X"54",X"3E",X"2D",X"06",X"01",X"21",X"88",X"D1",X"CD",X"15",X"54",X"3E",X"29",
		X"06",X"01",X"21",X"88",X"D2",X"CD",X"15",X"54",X"21",X"F8",X"D0",X"CD",X"28",X"54",X"21",X"F8",
		X"D2",X"CD",X"28",X"54",X"21",X"E8",X"D0",X"CD",X"28",X"54",X"CD",X"3C",X"54",X"CD",X"47",X"5E",
		X"CD",X"9C",X"5E",X"DD",X"E5",X"FD",X"E5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"FD",X"E1",X"DD",
		X"E1",X"DD",X"35",X"01",X"20",X"12",X"DD",X"36",X"01",X"4E",X"CD",X"CA",X"53",X"21",X"00",X"60",
		X"CB",X"E6",X"DD",X"35",X"00",X"CA",X"29",X"53",X"3A",X"65",X"60",X"A7",X"20",X"05",X"3A",X"00",
		X"90",X"18",X"03",X"3A",X"01",X"90",X"2F",X"E6",X"0F",X"28",X"C5",X"1F",X"38",X"68",X"1F",X"38",
		X"44",X"1F",X"38",X"21",X"FD",X"36",X"00",X"82",X"FD",X"7E",X"02",X"FE",X"D6",X"D2",X"E0",X"51",
		X"FD",X"4E",X"01",X"21",X"BD",X"53",X"CD",X"9F",X"53",X"D2",X"E0",X"51",X"FD",X"71",X"01",X"FD",
		X"34",X"02",X"C3",X"E0",X"51",X"FD",X"36",X"00",X"42",X"FD",X"7E",X"01",X"FE",X"A8",X"D2",X"E0",
		X"51",X"FD",X"4E",X"02",X"21",X"B1",X"53",X"CD",X"9F",X"53",X"D2",X"E0",X"51",X"FD",X"71",X"02",
		X"FD",X"34",X"01",X"18",X"3F",X"FD",X"36",X"00",X"22",X"FD",X"7E",X"02",X"FE",X"37",X"DA",X"E0",
		X"51",X"FD",X"4E",X"01",X"21",X"BD",X"53",X"CD",X"9F",X"53",X"D2",X"E0",X"51",X"FD",X"71",X"01",
		X"FD",X"35",X"02",X"C3",X"E0",X"51",X"FD",X"36",X"00",X"12",X"FD",X"7E",X"01",X"FE",X"09",X"DA",
		X"E0",X"51",X"FD",X"4E",X"02",X"21",X"B1",X"53",X"CD",X"9F",X"53",X"D2",X"E0",X"51",X"FD",X"71",
		X"02",X"FD",X"35",X"01",X"78",X"D6",X"02",X"DA",X"E0",X"51",X"FE",X"09",X"D2",X"E0",X"51",X"47",
		X"87",X"87",X"80",X"57",X"FD",X"4E",X"01",X"21",X"C4",X"53",X"CD",X"9F",X"53",X"A7",X"C2",X"E0",
		X"51",X"78",X"3D",X"82",X"5F",X"16",X"00",X"21",X"94",X"54",X"19",X"7E",X"A7",X"20",X"07",X"21",
		X"00",X"60",X"CB",X"FE",X"18",X"53",X"FE",X"80",X"20",X"1F",X"21",X"01",X"60",X"CB",X"CE",X"DD",
		X"7E",X"03",X"A7",X"CA",X"E0",X"51",X"DD",X"35",X"03",X"21",X"10",X"68",X"11",X"11",X"68",X"01",
		X"09",X"00",X"ED",X"B8",X"EB",X"36",X"FF",X"18",X"21",X"47",X"21",X"00",X"60",X"CB",X"C6",X"DD",
		X"7E",X"03",X"DD",X"BE",X"02",X"D2",X"E0",X"51",X"DD",X"34",X"03",X"C5",X"21",X"09",X"68",X"11",
		X"08",X"68",X"01",X"09",X"00",X"ED",X"B0",X"EB",X"C1",X"70",X"01",X"07",X"0A",X"11",X"08",X"68",
		X"21",X"7D",X"D1",X"CD",X"3F",X"5D",X"C3",X"E0",X"51",X"21",X"08",X"68",X"06",X"0A",X"3E",X"FF",
		X"BE",X"20",X"0E",X"23",X"10",X"FA",X"21",X"8A",X"54",X"11",X"08",X"68",X"01",X"0A",X"00",X"ED",
		X"B0",X"11",X"8D",X"60",X"DD",X"7E",X"04",X"D6",X"08",X"30",X"0D",X"ED",X"44",X"47",X"87",X"80",
		X"4F",X"06",X"00",X"21",X"8A",X"60",X"ED",X"B8",X"21",X"07",X"68",X"01",X"03",X"00",X"ED",X"B8",
		X"11",X"EB",X"D3",X"DD",X"7E",X"04",X"D6",X"08",X"30",X"0F",X"ED",X"44",X"87",X"87",X"47",X"87",
		X"80",X"4F",X"06",X"00",X"21",X"DF",X"D3",X"ED",X"B8",X"3E",X"FF",X"12",X"1B",X"21",X"11",X"68",
		X"01",X"0A",X"00",X"ED",X"B8",X"12",X"AF",X"32",X"26",X"60",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",
		X"21",X"80",X"D0",X"01",X"18",X"20",X"CD",X"52",X"5D",X"C9",X"00",X"00",X"00",X"00",X"C9",X"46",
		X"23",X"7E",X"91",X"30",X"02",X"ED",X"44",X"FE",X"07",X"38",X"04",X"23",X"10",X"F3",X"C9",X"4E",
		X"C9",X"0B",X"36",X"46",X"56",X"66",X"76",X"86",X"96",X"A6",X"B6",X"C6",X"D6",X"06",X"08",X"28",
		X"48",X"68",X"88",X"A8",X"05",X"1B",X"3B",X"5B",X"7B",X"9B",X"DD",X"7E",X"00",X"FE",X"0C",X"38",
		X"2C",X"FE",X"23",X"38",X"1F",X"FE",X"3A",X"38",X"14",X"FE",X"51",X"38",X"09",X"D6",X"5C",X"ED",
		X"44",X"11",X"1C",X"D6",X"18",X"1E",X"D6",X"3A",X"11",X"65",X"D7",X"18",X"21",X"D6",X"23",X"11",
		X"85",X"D4",X"18",X"10",X"D6",X"22",X"ED",X"44",X"11",X"86",X"D4",X"18",X"11",X"D6",X"0B",X"ED",
		X"44",X"11",X"BC",X"D4",X"6F",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"18",X"03",X"6F",X"26",
		X"00",X"19",X"36",X"05",X"C9",X"11",X"00",X"04",X"C5",X"E5",X"77",X"19",X"36",X"05",X"E1",X"01",
		X"80",X"00",X"09",X"C1",X"3C",X"10",X"F1",X"C9",X"01",X"20",X"00",X"11",X"00",X"04",X"E5",X"36",
		X"0C",X"19",X"36",X"06",X"E1",X"09",X"36",X"15",X"19",X"36",X"06",X"C9",X"3E",X"57",X"32",X"E8",
		X"D2",X"3C",X"32",X"08",X"D3",X"3E",X"07",X"32",X"E8",X"D6",X"32",X"08",X"D7",X"C9",X"DE",X"D0",
		X"06",X"07",X"22",X"18",X"1E",X"FF",X"10",X"0E",X"1D",X"5E",X"D2",X"06",X"08",X"11",X"12",X"FF",
		X"1C",X"0C",X"18",X"1B",X"0E",X"DD",X"D2",X"07",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1D",
		X"18",X"19",X"02",X"17",X"0D",X"03",X"1B",X"0D",X"04",X"1D",X"11",X"05",X"1D",X"11",X"06",X"1D",
		X"11",X"07",X"1D",X"11",X"08",X"1D",X"11",X"09",X"1D",X"11",X"FF",X"FF",X"15",X"0A",X"0D",X"22",
		X"FF",X"0B",X"1E",X"10",X"80",X"0C",X"0B",X"0A",X"80",X"11",X"10",X"0F",X"0E",X"0D",X"16",X"15",
		X"14",X"13",X"12",X"1B",X"1A",X"19",X"18",X"17",X"20",X"1F",X"1E",X"1D",X"1C",X"02",X"01",X"23",
		X"22",X"21",X"07",X"06",X"05",X"04",X"03",X"24",X"28",X"27",X"09",X"08",X"00",X"29",X"FF",X"2D",
		X"80",X"F5",X"C5",X"D5",X"E5",X"FD",X"E5",X"CD",X"9C",X"5D",X"21",X"C3",X"55",X"CD",X"1B",X"57",
		X"3E",X"C1",X"0E",X"08",X"21",X"D8",X"55",X"06",X"05",X"C5",X"5E",X"23",X"56",X"23",X"46",X"23",
		X"E5",X"EB",X"CD",X"C9",X"55",X"E1",X"C1",X"10",X"F0",X"3E",X"C0",X"21",X"D8",X"55",X"06",X"05",
		X"C5",X"5E",X"23",X"56",X"23",X"46",X"23",X"E5",X"EB",X"2B",X"CD",X"C9",X"55",X"E1",X"C1",X"10",
		X"EF",X"21",X"E7",X"55",X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",X"EB",
		X"CD",X"36",X"5D",X"FD",X"21",X"12",X"68",X"FD",X"36",X"00",X"22",X"FD",X"36",X"01",X"58",X"FD",
		X"36",X"02",X"D6",X"FD",X"36",X"03",X"10",X"FD",X"E5",X"CD",X"AE",X"5E",X"CD",X"C7",X"1F",X"CD",
		X"8F",X"17",X"FD",X"E1",X"FD",X"35",X"03",X"20",X"EE",X"21",X"B4",X"55",X"FD",X"74",X"04",X"FD",
		X"75",X"05",X"21",X"01",X"60",X"CB",X"D6",X"FD",X"66",X"04",X"FD",X"6E",X"05",X"7E",X"A7",X"28",
		X"41",X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"03",X"23",X"FD",X"74",X"04",X"FD",X"75",X"05",
		X"FD",X"7E",X"00",X"17",X"38",X"15",X"17",X"38",X"0D",X"17",X"38",X"05",X"FD",X"35",X"01",X"18",
		X"0D",X"FD",X"35",X"02",X"18",X"08",X"FD",X"34",X"01",X"18",X"03",X"FD",X"34",X"02",X"FD",X"E5",
		X"CD",X"AE",X"5E",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"FD",X"E1",X"FD",X"35",X"03",X"20",X"D0",
		X"18",X"B5",X"21",X"3F",X"60",X"36",X"00",X"FD",X"36",X"03",X"10",X"FD",X"E5",X"CD",X"C7",X"1F",
		X"CD",X"8F",X"17",X"FD",X"E1",X"FD",X"35",X"03",X"20",X"F1",X"CD",X"9C",X"5D",X"FD",X"E1",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"22",X"40",X"12",X"10",X"22",X"20",X"42",X"20",X"82",X"20",X"12",X"60",
		X"22",X"78",X"00",X"17",X"D1",X"03",X"10",X"C2",X"0B",X"11",X"00",X"04",X"E5",X"77",X"19",X"71",
		X"E1",X"11",X"20",X"00",X"19",X"10",X"F2",X"C9",X"F5",X"D0",X"07",X"55",X"D2",X"07",X"F1",X"D1",
		X"02",X"EF",X"D0",X"05",X"8F",X"D2",X"05",X"0C",X"D1",X"02",X"10",X"0C",X"18",X"17",X"10",X"1B",
		X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"28",X"AA",X"D1",X"02",X"07",X"22",
		X"18",X"1E",X"FF",X"20",X"12",X"17",X"28",X"D1",X"06",X"05",X"0E",X"21",X"1D",X"1B",X"0A",X"E8",
		X"D1",X"02",X"08",X"15",X"0A",X"0D",X"22",X"FF",X"0B",X"1E",X"10",X"F5",X"08",X"F5",X"C5",X"D5",
		X"E5",X"FD",X"E5",X"CD",X"9C",X"5D",X"FD",X"21",X"12",X"68",X"3A",X"27",X"60",X"FD",X"77",X"01",
		X"3A",X"28",X"60",X"FD",X"77",X"02",X"21",X"67",X"57",X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",
		X"06",X"10",X"CD",X"10",X"57",X"21",X"01",X"60",X"CB",X"DE",X"21",X"43",X"57",X"CD",X"1B",X"57",
		X"21",X"49",X"57",X"CD",X"1B",X"57",X"06",X"18",X"CD",X"10",X"57",X"21",X"4F",X"57",X"CD",X"1B",
		X"57",X"21",X"55",X"57",X"CD",X"1B",X"57",X"21",X"5B",X"57",X"CD",X"1B",X"57",X"21",X"73",X"57",
		X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",X"06",X"48",X"CD",X"10",X"57",X"21",X"61",X"57",X"CD",
		X"1B",X"57",X"3E",X"0A",X"32",X"09",X"D6",X"32",X"29",X"D6",X"06",X"30",X"CD",X"10",X"57",X"21",
		X"91",X"57",X"06",X"06",X"C5",X"CD",X"36",X"5D",X"C1",X"EB",X"10",X"F8",X"06",X"30",X"CD",X"10",
		X"57",X"FD",X"21",X"12",X"68",X"FD",X"7E",X"01",X"FE",X"0F",X"28",X"1D",X"38",X"09",X"FD",X"36",
		X"00",X"12",X"FD",X"35",X"01",X"18",X"07",X"FD",X"36",X"00",X"42",X"FD",X"34",X"01",X"CD",X"9C",
		X"5E",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"18",X"D8",X"FD",X"21",X"12",X"68",X"FD",X"7E",X"02",
		X"FE",X"CF",X"28",X"1D",X"38",X"09",X"FD",X"36",X"00",X"22",X"FD",X"35",X"02",X"18",X"07",X"FD",
		X"36",X"00",X"82",X"FD",X"34",X"02",X"CD",X"9C",X"5E",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"18",
		X"D8",X"01",X"02",X"02",X"21",X"D9",X"D0",X"CD",X"52",X"5D",X"AF",X"32",X"26",X"60",X"01",X"15",
		X"15",X"21",X"C6",X"D0",X"CD",X"52",X"5D",X"FD",X"E1",X"E1",X"D1",X"C1",X"F1",X"08",X"F1",X"C9",
		X"C5",X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"C1",X"10",X"F6",X"C9",X"5E",X"23",X"56",X"23",X"46",
		X"23",X"4E",X"23",X"7E",X"23",X"08",X"7E",X"08",X"EB",X"C5",X"E5",X"11",X"00",X"04",X"E5",X"77",
		X"19",X"08",X"77",X"08",X"3C",X"E1",X"23",X"10",X"F5",X"E1",X"11",X"20",X"00",X"19",X"C1",X"0D",
		X"20",X"E7",X"C9",X"C6",X"D0",X"08",X"06",X"10",X"0C",X"86",X"D2",X"08",X"06",X"90",X"0C",X"CC",
		X"D1",X"08",X"04",X"40",X"0A",X"88",X"D1",X"08",X"02",X"60",X"0A",X"48",X"D2",X"08",X"02",X"70",
		X"0A",X"C8",X"D1",X"04",X"04",X"00",X"0B",X"D9",X"D0",X"02",X"02",X"E9",X"E6",X"DA",X"D0",X"02",
		X"02",X"E8",X"E7",X"46",X"D1",X"0A",X"0C",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"88",X"67",X"D1",X"0A",X"0A",X"82",X"83",X"84",X"81",X"81",X"81",X"81",X"85",X"86",
		X"87",X"71",X"D1",X"07",X"01",X"29",X"93",X"D1",X"07",X"01",X"29",X"D4",X"D1",X"07",X"01",X"29",
		X"34",X"D2",X"07",X"01",X"29",X"73",X"D2",X"07",X"01",X"29",X"91",X"D2",X"07",X"01",X"29",X"21",
		X"00",X"B0",X"36",X"9F",X"36",X"BF",X"36",X"DF",X"36",X"FF",X"21",X"00",X"C0",X"36",X"9F",X"36",
		X"BF",X"36",X"DF",X"36",X"FF",X"21",X"00",X"D0",X"36",X"FF",X"23",X"7C",X"FE",X"D4",X"38",X"F8",
		X"36",X"00",X"23",X"7C",X"FE",X"D8",X"38",X"F8",X"0E",X"40",X"11",X"20",X"00",X"21",X"00",X"70",
		X"06",X"20",X"36",X"00",X"19",X"10",X"FB",X"0D",X"20",X"F3",X"21",X"00",X"00",X"AF",X"06",X"60",
		X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"A7",X"00",X"00",X"D9",X"47",X"D9",X"D9",X"0E",X"00",
		X"D9",X"1E",X"FF",X"21",X"00",X"60",X"16",X"10",X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",X"77",
		X"23",X"10",X"FA",X"3D",X"0D",X"20",X"F4",X"3D",X"15",X"20",X"EE",X"21",X"00",X"60",X"16",X"10",
		X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",X"BE",X"28",X"04",X"D9",X"0E",X"FF",X"D9",X"23",X"10",
		X"F4",X"3D",X"0D",X"20",X"EE",X"3D",X"15",X"20",X"E8",X"7B",X"D6",X"0F",X"5F",X"30",X"C4",X"3E",
		X"1B",X"32",X"92",X"D1",X"32",X"8F",X"D1",X"3E",X"18",X"32",X"B2",X"D1",X"3E",X"0A",X"32",X"AF",
		X"D1",X"3E",X"16",X"32",X"D2",X"D1",X"32",X"CF",X"D1",X"D9",X"78",X"A7",X"20",X"0C",X"3E",X"18",
		X"32",X"12",X"D2",X"3E",X"14",X"32",X"32",X"D2",X"18",X"1C",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",
		X"32",X"92",X"D2",X"78",X"E6",X"0F",X"32",X"B2",X"D2",X"3E",X"0E",X"32",X"12",X"D2",X"3E",X"1B",
		X"32",X"32",X"D2",X"32",X"52",X"D2",X"79",X"A7",X"20",X"0C",X"3E",X"18",X"32",X"0F",X"D2",X"3E",
		X"14",X"32",X"2F",X"D2",X"18",X"0D",X"3E",X"0E",X"32",X"0F",X"D2",X"3E",X"1B",X"32",X"2F",X"D2",
		X"32",X"4F",X"D2",X"78",X"B1",X"D9",X"11",X"03",X"00",X"28",X"03",X"11",X"12",X"00",X"01",X"00",
		X"00",X"0B",X"78",X"B1",X"20",X"FB",X"1B",X"7A",X"B3",X"20",X"F6",X"C3",X"00",X"01",X"A2",X"CD",
		X"9C",X"5D",X"CD",X"E5",X"1B",X"21",X"FF",X"5A",X"06",X"0D",X"C5",X"CD",X"36",X"5D",X"EB",X"C1",
		X"10",X"F8",X"CD",X"47",X"5E",X"DD",X"21",X"1A",X"68",X"DD",X"36",X"00",X"FF",X"3A",X"DF",X"5A",
		X"DD",X"77",X"01",X"21",X"E0",X"5A",X"DD",X"74",X"02",X"DD",X"75",X"03",X"DD",X"36",X"04",X"07",
		X"DD",X"36",X"05",X"1E",X"DD",X"36",X"06",X"00",X"FD",X"21",X"12",X"68",X"FD",X"36",X"00",X"42",
		X"FD",X"36",X"01",X"08",X"FD",X"36",X"02",X"B7",X"CD",X"9C",X"5E",X"DD",X"E5",X"FD",X"E5",X"CD",
		X"C7",X"1F",X"CD",X"8F",X"17",X"FD",X"E1",X"DD",X"E1",X"DD",X"35",X"05",X"20",X"07",X"DD",X"36",
		X"05",X"1E",X"CD",X"93",X"5A",X"DD",X"7E",X"00",X"A7",X"28",X"08",X"DD",X"35",X"01",X"CC",X"7A",
		X"5A",X"18",X"D5",X"FD",X"34",X"01",X"DD",X"35",X"01",X"20",X"CD",X"CD",X"44",X"5A",X"DD",X"7E",
		X"06",X"FE",X"0F",X"30",X"28",X"CD",X"B8",X"59",X"CD",X"7A",X"5A",X"DD",X"34",X"06",X"DD",X"7E",
		X"06",X"FE",X"0C",X"28",X"0E",X"FE",X"05",X"20",X"AF",X"FD",X"36",X"01",X"08",X"FD",X"36",X"02",
		X"9F",X"18",X"A5",X"FD",X"36",X"01",X"08",X"FD",X"36",X"02",X"87",X"18",X"9B",X"3E",X"81",X"32",
		X"26",X"60",X"21",X"9A",X"59",X"0E",X"0F",X"06",X"1E",X"5E",X"23",X"56",X"23",X"ED",X"53",X"29",
		X"60",X"C5",X"E5",X"CD",X"10",X"57",X"E1",X"C1",X"06",X"05",X"0D",X"20",X"EC",X"06",X"3C",X"CD",
		X"10",X"57",X"AF",X"32",X"26",X"60",X"C3",X"F0",X"5E",X"C9",X"E4",X"00",X"E8",X"00",X"EC",X"00",
		X"F0",X"00",X"F4",X"00",X"F8",X"00",X"FC",X"00",X"FC",X"09",X"48",X"19",X"4C",X"19",X"50",X"19",
		X"54",X"19",X"58",X"19",X"5C",X"19",X"60",X"19",X"DD",X"7E",X"06",X"FE",X"0C",X"30",X"37",X"FE",
		X"05",X"30",X"17",X"CD",X"20",X"5A",X"11",X"DD",X"D5",X"19",X"36",X"06",X"FE",X"04",X"C0",X"21",
		X"2C",X"5A",X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",X"C9",X"D6",X"05",X"CD",X"20",X"5A",X"11",
		X"BD",X"D4",X"19",X"36",X"07",X"DD",X"7E",X"06",X"FE",X"0B",X"C0",X"21",X"38",X"5A",X"CD",X"36",
		X"5D",X"EB",X"CD",X"36",X"5D",X"C9",X"D6",X"0C",X"87",X"CD",X"20",X"5A",X"11",X"BD",X"D6",X"19",
		X"36",X"05",X"11",X"20",X"00",X"19",X"36",X"05",X"0F",X"5F",X"16",X"00",X"21",X"29",X"5A",X"19",
		X"3E",X"56",X"32",X"ED",X"D2",X"32",X"EA",X"D2",X"7E",X"32",X"0D",X"D3",X"32",X"0A",X"D3",X"C9",
		X"6F",X"26",X"00",X"29",X"29",X"29",X"29",X"29",X"C9",X"02",X"03",X"05",X"17",X"D3",X"01",X"02",
		X"E3",X"E4",X"16",X"D3",X"01",X"02",X"E1",X"E2",X"14",X"D3",X"02",X"02",X"E8",X"E7",X"13",X"D3",
		X"02",X"02",X"E9",X"E6",X"DD",X"7E",X"06",X"87",X"5F",X"16",X"00",X"21",X"5A",X"5A",X"19",X"5E",
		X"23",X"56",X"EB",X"01",X"02",X"02",X"CD",X"52",X"5D",X"C9",X"36",X"D1",X"76",X"D1",X"B6",X"D1",
		X"F6",X"D1",X"36",X"D2",X"33",X"D1",X"73",X"D1",X"B3",X"D1",X"F3",X"D1",X"33",X"D2",X"73",X"D2",
		X"B3",X"D2",X"30",X"D1",X"B0",X"D1",X"30",X"D2",X"10",X"D3",X"DD",X"7E",X"00",X"2F",X"DD",X"77",
		X"00",X"DD",X"66",X"02",X"DD",X"6E",X"03",X"7E",X"DD",X"77",X"01",X"23",X"DD",X"74",X"02",X"DD",
		X"75",X"03",X"C9",X"DD",X"7E",X"04",X"3D",X"FE",X"05",X"30",X"02",X"3E",X"07",X"DD",X"77",X"04",
		X"21",X"37",X"D5",X"06",X"0A",X"CD",X"CA",X"5A",X"2B",X"06",X"0E",X"CD",X"CA",X"5A",X"2B",X"06",
		X"0A",X"CD",X"CA",X"5A",X"21",X"2B",X"D5",X"06",X"02",X"CD",X"CA",X"5A",X"D6",X"05",X"5F",X"16",
		X"00",X"21",X"DC",X"5A",X"19",X"7E",X"32",X"8A",X"D1",X"C9",X"0E",X"02",X"11",X"20",X"00",X"C5",
		X"E5",X"77",X"19",X"10",X"FC",X"E1",X"2B",X"C1",X"0D",X"20",X"F4",X"C9",X"01",X"03",X"08",X"68",
		X"20",X"4A",X"10",X"4A",X"10",X"4A",X"10",X"4A",X"10",X"1C",X"20",X"4A",X"10",X"4A",X"10",X"4A",
		X"10",X"4A",X"10",X"4A",X"10",X"4A",X"10",X"1C",X"20",X"3A",X"20",X"3A",X"20",X"3A",X"38",X"79",
		X"D1",X"02",X"0B",X"12",X"17",X"1C",X"1D",X"1B",X"1E",X"0C",X"1D",X"12",X"18",X"17",X"37",X"D1",
		X"07",X"0A",X"F1",X"65",X"F4",X"6D",X"F5",X"6F",X"F1",X"67",X"F1",X"67",X"36",X"D1",X"07",X"0A",
		X"95",X"5B",X"9D",X"5F",X"9F",X"60",X"93",X"61",X"9B",X"5E",X"34",X"D1",X"07",X"0E",X"F1",X"65",
		X"F1",X"67",X"F1",X"65",X"F1",X"65",X"F2",X"69",X"F1",X"67",X"F3",X"6B",X"33",X"D1",X"07",X"0E",
		X"91",X"59",X"93",X"5A",X"95",X"5B",X"97",X"5C",X"99",X"5D",X"9B",X"5E",X"97",X"5C",X"31",X"D1",
		X"07",X"0A",X"EF",X"71",X"FF",X"FF",X"EF",X"71",X"FF",X"FF",X"EF",X"71",X"30",X"D1",X"07",X"0A",
		X"A1",X"62",X"FF",X"FF",X"A1",X"62",X"FF",X"FF",X"A1",X"62",X"11",X"D3",X"06",X"02",X"F0",X"73",
		X"10",X"D3",X"06",X"02",X"A3",X"63",X"4D",X"D1",X"02",X"0F",X"E5",X"FF",X"FF",X"01",X"00",X"FF",
		X"19",X"18",X"12",X"17",X"1D",X"1C",X"FF",X"FF",X"FF",X"2B",X"D1",X"07",X"02",X"F4",X"6D",X"2A",
		X"D1",X"07",X"02",X"9D",X"5F",X"8A",X"D1",X"02",X"0D",X"08",X"00",X"00",X"FF",X"19",X"18",X"12",
		X"17",X"1D",X"1C",X"FF",X"FF",X"FF",X"C3",X"00",X"5F",X"11",X"1C",X"60",X"01",X"32",X"00",X"ED",
		X"B0",X"21",X"56",X"5C",X"CD",X"36",X"5D",X"3A",X"03",X"90",X"E6",X"0F",X"F5",X"21",X"26",X"D1",
		X"CD",X"41",X"5C",X"F1",X"47",X"3E",X"06",X"32",X"26",X"D5",X"32",X"26",X"D6",X"3A",X"03",X"90",
		X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"B8",X"C8",X"21",X"23",X"D1",X"CD",X"41",X"5C",X"3E",X"06",
		X"32",X"23",X"D5",X"32",X"23",X"D6",X"21",X"1B",X"5D",X"CD",X"36",X"5D",X"EB",X"CD",X"36",X"5D",
		X"C9",X"F5",X"C5",X"06",X"1F",X"CD",X"10",X"57",X"C1",X"F1",X"C9",X"21",X"1C",X"60",X"36",X"00",
		X"11",X"1D",X"60",X"01",X"31",X"00",X"ED",X"B0",X"CD",X"C7",X"1F",X"C3",X"10",X"5F",X"C9",X"42",
		X"17",X"AF",X"30",X"02",X"82",X"3F",X"DF",X"78",X"05",X"82",X"5F",X"A7",X"60",X"04",X"12",X"97",
		X"CF",X"18",X"01",X"42",X"10",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E5",X"87",X"5F",X"16",X"00",X"21",X"65",X"5C",X"19",X"5E",X"23",X"56",X"E1",X"06",X"0F",
		X"0E",X"02",X"CD",X"3F",X"5D",X"C9",X"69",X"D1",X"00",X"0B",X"12",X"17",X"1C",X"0E",X"1B",X"1D",
		X"FF",X"0C",X"18",X"12",X"17",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",X"5C",X"85",
		X"5C",X"0C",X"5D",X"FD",X"5C",X"EE",X"5C",X"DF",X"5C",X"D0",X"5C",X"C1",X"5C",X"B2",X"5C",X"A3",
		X"5C",X"94",X"5C",X"85",X"5C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"01",X"FF",X"19",
		X"15",X"0A",X"22",X"FF",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"02",X"FF",X"19",X"15",
		X"0A",X"22",X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"03",X"FF",X"19",X"15",X"0A",
		X"22",X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"04",X"FF",X"19",X"15",X"0A",X"22",
		X"1C",X"01",X"FF",X"0C",X"18",X"12",X"17",X"FF",X"FF",X"05",X"FF",X"19",X"15",X"0A",X"22",X"1C",
		X"02",X"FF",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"02",
		X"FF",X"0C",X"18",X"12",X"17",X"1C",X"FF",X"03",X"FF",X"19",X"15",X"0A",X"22",X"1C",X"03",X"FF",
		X"0C",X"18",X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"03",X"FF",X"0C",
		X"18",X"12",X"17",X"1C",X"FF",X"02",X"FF",X"19",X"15",X"0A",X"22",X"1C",X"04",X"FF",X"0C",X"18",
		X"12",X"17",X"1C",X"FF",X"01",X"FF",X"19",X"15",X"0A",X"22",X"FF",X"E7",X"D0",X"01",X"05",X"1B",
		X"12",X"10",X"11",X"1D",X"E4",X"D0",X"01",X"04",X"15",X"0E",X"0F",X"1D",X"06",X"03",X"1A",X"BE",
		X"C0",X"13",X"23",X"10",X"F9",X"C9",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"EB",X"D5",
		X"E5",X"1A",X"77",X"11",X"00",X"04",X"19",X"71",X"E1",X"11",X"20",X"00",X"19",X"D1",X"13",X"10",
		X"EE",X"C9",X"D5",X"11",X"00",X"04",X"C5",X"E5",X"E5",X"36",X"FF",X"19",X"36",X"00",X"E1",X"23",
		X"10",X"F6",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",X"20",X"EB",X"D1",X"C9",X"11",X"DD",X"D2",
		X"21",X"05",X"68",X"AF",X"06",X"06",X"ED",X"6F",X"28",X"09",X"F6",X"80",X"F5",X"E6",X"0F",X"C6",
		X"00",X"12",X"F1",X"E5",X"21",X"20",X"00",X"19",X"EB",X"E1",X"CB",X"40",X"28",X"05",X"ED",X"6F",
		X"23",X"18",X"06",X"CB",X"48",X"20",X"02",X"F6",X"80",X"10",X"DB",X"C9",X"01",X"18",X"18",X"21",
		X"85",X"D0",X"CD",X"52",X"5D",X"21",X"1C",X"60",X"11",X"05",X"00",X"36",X"00",X"19",X"36",X"00",
		X"19",X"06",X"07",X"19",X"36",X"00",X"10",X"FB",X"CD",X"BC",X"5D",X"C9",X"0E",X"06",X"3E",X"4E",
		X"32",X"9C",X"D0",X"79",X"32",X"9C",X"D4",X"3E",X"4F",X"32",X"7C",X"D3",X"79",X"32",X"7C",X"D7",
		X"3E",X"51",X"32",X"85",X"D0",X"79",X"32",X"85",X"D4",X"3E",X"50",X"32",X"65",X"D3",X"79",X"32",
		X"65",X"D7",X"3E",X"52",X"06",X"16",X"21",X"BC",X"D0",X"CD",X"2A",X"5E",X"3E",X"54",X"06",X"16",
		X"21",X"A5",X"D0",X"CD",X"2A",X"5E",X"3E",X"55",X"06",X"16",X"21",X"86",X"D0",X"CD",X"3B",X"5E",
		X"3E",X"53",X"06",X"16",X"21",X"66",X"D3",X"CD",X"3B",X"5E",X"0E",X"00",X"3E",X"30",X"32",X"BB",
		X"D0",X"79",X"32",X"BB",X"D4",X"3E",X"31",X"06",X"15",X"21",X"DB",X"D0",X"CD",X"2A",X"5E",X"3E",
		X"32",X"06",X"15",X"21",X"A6",X"D0",X"CD",X"3B",X"5E",X"C9",X"11",X"00",X"04",X"C5",X"E5",X"77",
		X"19",X"71",X"E1",X"01",X"20",X"00",X"09",X"C1",X"10",X"F3",X"C9",X"11",X"00",X"04",X"E5",X"77",
		X"19",X"71",X"E1",X"23",X"10",X"F8",X"C9",X"DD",X"E5",X"FD",X"E5",X"CD",X"D1",X"1D",X"CD",X"8B",
		X"1E",X"06",X"06",X"3E",X"05",X"21",X"A1",X"D5",X"CD",X"7D",X"1E",X"CD",X"E0",X"1E",X"CD",X"26",
		X"28",X"06",X"05",X"3E",X"01",X"21",X"E1",X"D4",X"CD",X"7D",X"1E",X"21",X"E1",X"D0",X"36",X"2A",
		X"19",X"CD",X"44",X"1F",X"DD",X"21",X"1C",X"60",X"DD",X"36",X"00",X"82",X"DD",X"36",X"01",X"08",
		X"DD",X"36",X"02",X"0F",X"CD",X"7F",X"1F",X"DD",X"77",X"03",X"DD",X"70",X"04",X"CD",X"C7",X"1F",
		X"CD",X"8F",X"17",X"DD",X"36",X"00",X"81",X"FD",X"E1",X"DD",X"E1",X"C9",X"11",X"26",X"60",X"21",
		X"12",X"68",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"36",X"00",X"23",X"36",X"00",X"C9",X"11",X"3F",
		X"60",X"18",X"EC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E6",X"02",X"CA",X"E3",X"5E",X"C3",X"78",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"A4",X"50",X"DA",X"E3",X"5E",X"C3",X"88",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"F6",X"50",X"CD",X"3E",X"25",X"CD",X"07",X"26",X"CD",X"B1",X"5B",X"00",X"00",X"00",X"C9",
		X"CD",X"C7",X"1F",X"CD",X"8F",X"17",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"32",X"65",X"60",X"21",X"0F",X"5C",X"C3",X"A9",X"5B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"8F",X"17",X"21",X"80",X"D0",X"01",X"18",X"20",X"CD",X"52",X"5D",X"C9",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
