library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_char_l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_char_l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"3C",X"66",X"42",X"42",X"42",X"66",X"3C",X"00",X"00",X"00",X"22",X"7E",X"02",X"00",X"00",
		X"00",X"26",X"6E",X"4A",X"4A",X"4A",X"7A",X"32",X"00",X"44",X"46",X"52",X"52",X"52",X"7E",X"6C",
		X"00",X"0C",X"1C",X"34",X"64",X"44",X"7E",X"04",X"00",X"74",X"56",X"52",X"52",X"52",X"5E",X"0C",
		X"00",X"3C",X"76",X"52",X"52",X"52",X"5E",X"0C",X"00",X"40",X"42",X"46",X"4C",X"58",X"70",X"60",
		X"00",X"2C",X"7E",X"52",X"52",X"52",X"7E",X"2C",X"00",X"30",X"7A",X"4A",X"4A",X"4A",X"6E",X"3C",
		X"00",X"1E",X"34",X"64",X"44",X"64",X"34",X"1E",X"00",X"7E",X"52",X"52",X"52",X"52",X"7E",X"2C",
		X"00",X"3C",X"66",X"42",X"42",X"42",X"66",X"24",X"00",X"7E",X"42",X"42",X"42",X"42",X"66",X"3C",
		X"00",X"7E",X"52",X"52",X"52",X"52",X"42",X"42",X"00",X"7E",X"50",X"50",X"50",X"50",X"40",X"40",
		X"00",X"3C",X"66",X"42",X"42",X"4A",X"6A",X"2E",X"00",X"7E",X"10",X"10",X"10",X"10",X"10",X"7E",
		X"00",X"00",X"00",X"42",X"7E",X"42",X"00",X"00",X"00",X"0C",X"06",X"02",X"02",X"02",X"06",X"7C",
		X"00",X"7E",X"06",X"0C",X"18",X"34",X"66",X"42",X"00",X"7E",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"7E",X"30",X"18",X"0C",X"18",X"30",X"7E",X"00",X"7E",X"60",X"30",X"18",X"0C",X"06",X"7E",
		X"00",X"3C",X"66",X"42",X"42",X"42",X"66",X"3C",X"00",X"7E",X"48",X"48",X"48",X"48",X"78",X"30",
		X"00",X"3C",X"66",X"42",X"4A",X"4C",X"66",X"3A",X"00",X"7E",X"48",X"48",X"48",X"4E",X"7A",X"32",
		X"00",X"24",X"76",X"52",X"5A",X"4A",X"6E",X"24",X"00",X"40",X"40",X"40",X"7E",X"40",X"40",X"40",
		X"00",X"7C",X"06",X"02",X"02",X"02",X"06",X"7C",X"00",X"70",X"1C",X"06",X"02",X"06",X"1C",X"70",
		X"00",X"7C",X"06",X"0C",X"18",X"0C",X"06",X"7C",X"00",X"42",X"66",X"2C",X"18",X"34",X"66",X"42",
		X"00",X"60",X"30",X"18",X"0E",X"18",X"30",X"60",X"00",X"42",X"46",X"4E",X"5A",X"72",X"62",X"42",
		X"00",X"6C",X"7E",X"52",X"42",X"16",X"1C",X"10",X"00",X"24",X"7E",X"24",X"24",X"24",X"7E",X"24",
		X"00",X"2E",X"6A",X"4E",X"42",X"42",X"66",X"3C",X"00",X"20",X"60",X"40",X"5A",X"50",X"70",X"20",
		X"00",X"00",X"00",X"00",X"7A",X"60",X"00",X"00",X"00",X"30",X"78",X"7C",X"3E",X"7C",X"78",X"30",
		X"00",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"00",X"00",X"18",X"3C",X"66",X"42",X"00",X"00",
		X"00",X"00",X"42",X"66",X"3C",X"18",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"00",X"7C",X"82",X"BA",X"AA",X"AA",X"82",X"7C",
		X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",
		X"FF",X"FF",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"00",X"C0",X"C0",X"C0",X"C0",X"C0",X"DF",X"DF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DF",X"DF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",
		X"00",X"00",X"30",X"38",X"1C",X"0E",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"0E",X"1C",X"38",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"0E",X"1C",X"38",X"30",
		X"C0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"14",X"08",X"14",X"22",X"00",X"7E",X"52",X"52",X"52",X"00",X"7E",X"30",
		X"18",X"0C",X"7E",X"00",X"7E",X"42",X"66",X"3C",X"58",X"58",X"10",X"F0",X"C0",X"00",X"00",X"00",
		X"78",X"78",X"70",X"F0",X"C0",X"00",X"00",X"00",X"58",X"58",X"D0",X"F0",X"C0",X"00",X"00",X"00",
		X"D8",X"D8",X"D0",X"F0",X"C0",X"00",X"00",X"00",X"18",X"D8",X"F0",X"F0",X"C0",X"00",X"00",X"00",
		X"B8",X"B8",X"10",X"F0",X"C0",X"00",X"00",X"00",X"78",X"38",X"90",X"F0",X"C0",X"00",X"00",X"00",
		X"18",X"F8",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"78",X"18",X"50",X"F0",X"C0",X"00",X"00",X"00",
		X"F8",X"F8",X"F0",X"F0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CD",X"CD",X"C5",X"C7",X"C1",X"C0",X"C0",X"C0",X"0D",X"0D",X"05",X"07",X"01",X"00",X"00",X"00",
		X"CD",X"CD",X"C4",X"C7",X"C1",X"C0",X"C0",X"C0",X"0D",X"0D",X"04",X"07",X"01",X"00",X"00",X"00",
		X"CC",X"CD",X"C7",X"C7",X"C1",X"C0",X"C0",X"C0",X"0C",X"0D",X"07",X"07",X"01",X"00",X"00",X"00",
		X"CF",X"CF",X"C7",X"C7",X"C1",X"C0",X"C0",X"C0",X"0F",X"0F",X"07",X"07",X"01",X"00",X"00",X"00",
		X"CF",X"CE",X"C4",X"C7",X"C1",X"C0",X"C0",X"C0",X"0F",X"0E",X"04",X"07",X"01",X"00",X"00",X"00",
		X"CC",X"CD",X"C5",X"C7",X"C1",X"C0",X"C0",X"C0",X"0C",X"0D",X"05",X"07",X"01",X"00",X"00",X"00",
		X"CF",X"CF",X"C7",X"C7",X"C1",X"C0",X"C0",X"C0",X"0F",X"0F",X"07",X"07",X"01",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C4",X"CD",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C4",X"CD",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"04",X"0D",X"C0",X"C0",X"00",X"00",X"01",X"07",X"04",X"0D",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C7",X"CD",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C7",X"CD",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"07",X"0D",X"C0",X"C0",X"00",X"00",X"01",X"07",X"07",X"0D",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C4",X"CF",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C4",X"CF",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"04",X"0F",X"C0",X"C0",X"00",X"00",X"01",X"07",X"04",X"0F",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C4",X"CE",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C4",X"CE",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"04",X"0E",X"C0",X"C0",X"00",X"00",X"01",X"07",X"04",X"0E",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C5",X"CD",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C5",X"CD",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"05",X"0D",X"C0",X"C0",X"00",X"00",X"01",X"07",X"05",X"0D",
		X"FF",X"FF",X"C0",X"C0",X"C1",X"C7",X"C7",X"CF",X"C0",X"C0",X"C0",X"C0",X"C1",X"C7",X"C7",X"CF",
		X"FF",X"FF",X"00",X"00",X"01",X"07",X"07",X"0F",X"C0",X"C0",X"00",X"00",X"01",X"07",X"07",X"0F",
		X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"50",X"58",X"00",X"00",X"00",X"00",X"C0",X"F0",X"50",X"58",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"10",X"78",X"00",X"00",X"00",X"00",X"C0",X"F0",X"10",X"78",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"10",X"58",X"00",X"00",X"00",X"00",X"C0",X"F0",X"10",X"58",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"10",X"D8",X"00",X"00",X"00",X"00",X"C0",X"F0",X"10",X"D8",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"F0",X"D8",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"D8",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"10",X"B8",X"00",X"00",X"00",X"00",X"C0",X"F0",X"10",X"B8",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"90",X"38",X"00",X"00",X"00",X"00",X"C0",X"F0",X"90",X"38",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F8",
		X"FF",X"FF",X"00",X"00",X"C0",X"F0",X"F0",X"F8",X"00",X"00",X"00",X"00",X"C0",X"F0",X"F0",X"F8",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"20",X"00",X"00",X"20",X"40",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"18",X"20",X"00",X"00",X"00",X"08",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"02",X"05",X"00",X"13",X"25",X"19",X"00",X"05",X"02",X"05",X"00",X"22",X"29",X"36",X"00",
		X"05",X"02",X"05",X"00",X"0E",X"12",X"3F",X"02",X"05",X"02",X"05",X"00",X"3A",X"29",X"26",X"00",
		X"05",X"02",X"05",X"00",X"1E",X"29",X"26",X"00",X"05",X"02",X"05",X"00",X"23",X"2C",X"30",X"00",
		X"05",X"02",X"05",X"00",X"16",X"29",X"16",X"00",X"00",X"00",X"00",X"40",X"00",X"90",X"C0",X"D8",
		X"98",X"00",X"00",X"00",X"E0",X"80",X"40",X"00",X"00",X"00",X"00",X"02",X"00",X"09",X"03",X"1B",
		X"19",X"00",X"00",X"00",X"07",X"01",X"02",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",X"00",
		X"07",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"C0",X"00",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"07",X"00",
		X"07",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",
		X"C0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"07",X"04",X"0D",
		X"00",X"00",X"00",X"00",X"01",X"07",X"07",X"0D",X"00",X"00",X"00",X"00",X"01",X"07",X"04",X"0F",
		X"00",X"00",X"00",X"00",X"01",X"07",X"04",X"0E",X"00",X"00",X"00",X"00",X"01",X"07",X"05",X"0D",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FE",X"00",X"00",X"00",X"00",X"30",X"30",X"3F",X"7F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",
		X"FE",X"00",X"FE",X"FE",X"FE",X"00",X"00",X"00",X"FF",X"F0",X"FF",X"7F",X"3F",X"00",X"C8",X"18",
		X"80",X"E1",X"80",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FE",X"FC",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"EF",X"FF",X"DF",X"AF",X"1F",X"AF",
		X"30",X"E1",X"C7",X"81",X"C0",X"E0",X"E0",X"C3",X"00",X"00",X"03",X"0F",X"3F",X"7F",X"7F",X"3F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DF",X"FF",X"EF",X"C3",X"00",X"00",X"00",X"00",
		X"80",X"C1",X"FF",X"3F",X"0F",X"00",X"00",X"00",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"13",X"3F",X"7F",X"CF",X"DF",X"7F",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"00",X"1E",X"3F",X"7F",X"FF",X"FF",X"00",X"00",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F1",X"FB",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"E3",X"F7",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"C0",X"E0",X"E0",X"F0",X"F0",X"E0",X"C7",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",
		X"7F",X"7F",X"3F",X"3F",X"1F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"07",X"03",X"1F",X"3F",X"3F",X"5F",X"FC",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"00",X"00",X"FF",X"FF",X"FF",X"FB",X"71",X"00",X"00",X"84",
		X"FF",X"FE",X"7C",X"00",X"00",X"02",X"3E",X"FF",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"7F",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"00",X"00",X"C0",X"C0",X"E0",X"F0",X"F0",X"F0",
		X"00",X"00",X"C1",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"37",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FE",X"FC",X"10",X"01",X"03",X"07",X"0F",X"1F",X"FF",X"FF",X"E0",X"C0",X"80",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EF",X"C7",X"02",X"10",X"F8",X"FF",X"F7",X"E3",X"01",X"10",X"FC",X"FE",X"FF",
		X"3F",X"07",X"03",X"00",X"02",X"0F",X"5F",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"1F",X"1F",X"0F",X"FF",X"07",X"03",X"00",X"00",X"C0",X"E0",X"E0",X"FF",X"E0",X"C0",X"00",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"67",X"03",
		X"FF",X"FF",X"FF",X"FF",X"1F",X"0E",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CF",X"9E",X"3C",X"7C",X"F8",X"F8",X"F8",X"F0",X"DF",X"EF",X"DF",X"EE",X"DC",X"F9",X"F3",X"E7",
		X"FF",X"3C",X"FF",X"3F",X"FF",X"3C",X"FF",X"3F",X"FE",X"62",X"6E",X"0E",X"6E",X"02",X"BE",X"7E",
		X"7F",X"D0",X"17",X"C7",X"D7",X"00",X"FF",X"FF",X"00",X"FF",X"38",X"83",X"BB",X"80",X"AF",X"9F",
		X"00",X"07",X"18",X"7B",X"FF",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"B0",X"CF",X"9F",X"3F",X"7F",X"F1",X"FD",X"8C",X"FF",
		X"FF",X"3F",X"FF",X"3E",X"FC",X"39",X"F3",X"E7",X"BE",X"FE",X"FE",X"7E",X"3E",X"1E",X"5E",X"FE",
		X"FF",X"FF",X"80",X"0F",X"7F",X"FF",X"FF",X"FF",X"AF",X"9F",X"AF",X"9F",X"AE",X"9C",X"AD",X"9F",
		X"03",X"00",X"01",X"03",X"06",X"0D",X"1B",X"F7",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"FF",
		X"B0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"9F",X"CF",
		X"E7",X"F3",X"39",X"FC",X"3E",X"FF",X"3F",X"FF",X"FE",X"5E",X"1E",X"3E",X"7E",X"FE",X"FE",X"BE",
		X"FF",X"FF",X"FF",X"7F",X"0F",X"80",X"FF",X"FF",X"AF",X"9D",X"AC",X"9E",X"AF",X"9F",X"AF",X"9F",
		X"F7",X"1B",X"0D",X"06",X"03",X"01",X"00",X"03",X"FF",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",
		X"F0",X"F8",X"F8",X"F8",X"7C",X"3C",X"9E",X"CF",X"E7",X"F3",X"F9",X"DC",X"EE",X"DF",X"EF",X"DF",
		X"3F",X"FF",X"3C",X"FF",X"3F",X"FF",X"3C",X"FF",X"7E",X"BE",X"06",X"6E",X"0E",X"6E",X"66",X"FE",
		X"FF",X"FF",X"00",X"D7",X"C7",X"17",X"D0",X"7F",X"AF",X"9F",X"80",X"BB",X"83",X"38",X"FF",X"00",
		X"00",X"03",X"00",X"FF",X"7B",X"18",X"07",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"F9",X"FA",X"39",X"3A",X"39",X"FA",X"F9",X"FF",X"FF",X"7F",X"FE",X"72",X"E2",X"7F",X"FF",
		X"FF",X"DA",X"B6",X"DA",X"B6",X"DA",X"B6",X"DA",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"FF",X"FF",
		X"FF",X"4F",X"D7",X"4F",X"D6",X"4F",X"D7",X"4F",X"FF",X"FD",X"FE",X"05",X"06",X"05",X"06",X"FD",
		X"FF",X"7F",X"BF",X"78",X"B0",X"70",X"B8",X"7F",X"07",X"1F",X"07",X"01",X"01",X"07",X"1F",X"FF",
		X"3A",X"39",X"3A",X"F9",X"FA",X"FF",X"00",X"00",X"62",X"F2",X"7E",X"FF",X"7F",X"FF",X"00",X"00",
		X"B6",X"DA",X"B6",X"DA",X"B6",X"FF",X"00",X"00",X"FF",X"01",X"01",X"01",X"FF",X"FF",X"FE",X"E0",
		X"D7",X"4F",X"D6",X"4F",X"DB",X"7B",X"F3",X"E7",X"FE",X"FD",X"06",X"05",X"06",X"05",X"FE",X"FD",
		X"BF",X"7F",X"B8",X"70",X"B0",X"78",X"BF",X"FF",X"1F",X"07",X"01",X"01",X"07",X"1F",X"07",X"01",
		X"00",X"00",X"FF",X"FA",X"F9",X"3A",X"39",X"3A",X"00",X"00",X"FF",X"7F",X"FF",X"7E",X"F2",X"62",
		X"00",X"00",X"FF",X"B6",X"DA",X"B6",X"DA",X"B6",X"E0",X"FE",X"FF",X"FF",X"01",X"01",X"01",X"FF",
		X"E7",X"F3",X"7B",X"DB",X"4F",X"D6",X"4F",X"D7",X"FD",X"FE",X"05",X"06",X"05",X"06",X"FD",X"FE",
		X"FF",X"BF",X"78",X"B0",X"70",X"B8",X"7F",X"BF",X"01",X"07",X"1F",X"07",X"01",X"01",X"07",X"1F",
		X"F9",X"FA",X"39",X"3A",X"39",X"FA",X"F9",X"FF",X"FF",X"7F",X"E2",X"72",X"FE",X"7F",X"FF",X"FF",
		X"DA",X"B6",X"DA",X"B6",X"DA",X"B6",X"DA",X"FF",X"FF",X"FF",X"01",X"01",X"01",X"FF",X"FF",X"FF",
		X"4F",X"D7",X"4F",X"D6",X"4F",X"D7",X"4F",X"FF",X"FD",X"06",X"05",X"06",X"05",X"FE",X"FD",X"FF",
		X"7F",X"B8",X"70",X"B0",X"78",X"BF",X"7F",X"FF",X"FF",X"1F",X"07",X"01",X"01",X"07",X"1F",X"07",
		X"03",X"03",X"0F",X"0F",X"3F",X"3F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"14",X"41",X"11",X"14",X"41",X"11",X"14",X"41",X"11",X"14",X"41",X"11",X"14",X"41",X"10",
		X"17",X"43",X"1F",X"0F",X"7F",X"3F",X"FF",X"FF",X"FF",X"FF",X"3F",X"7F",X"0F",X"1F",X"43",X"17",
		X"10",X"41",X"14",X"11",X"41",X"14",X"11",X"41",X"14",X"11",X"41",X"14",X"11",X"41",X"14",X"01",
		X"FF",X"FF",X"3F",X"3F",X"0F",X"0F",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"07",X"FF",X"0F",X"1F",X"1F",X"1F",X"00",X"C0",X"E0",X"FF",X"E0",X"E0",X"C0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"03",X"67",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"0E",X"1F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"0F",X"07",X"03",X"01",X"10",X"FC",X"FE",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FF",X"FF",
		X"F8",X"10",X"02",X"C7",X"EF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"10",X"01",X"E3",X"F7",X"FF",
		X"FF",X"5F",X"0F",X"02",X"00",X"03",X"07",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"7F",X"7F",X"F0",X"F0",X"F0",X"E0",X"C0",X"C0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",
		X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"37",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"5F",X"3F",X"3F",X"1F",X"03",X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",X"FC",
		X"00",X"00",X"7C",X"FF",X"FF",X"FF",X"FF",X"FF",X"84",X"00",X"00",X"71",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"3E",X"02",X"00",X"00",X"7C",X"FE",X"FF",X"0B",X"00",X"00",X"00",X"00",X"00",X"03",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"3F",X"FF",X"C7",X"E0",X"F0",X"F0",X"E0",X"E0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"03",X"07",X"1F",X"3F",X"3F",X"7F",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"DF",X"CF",X"7F",X"3F",X"13",X"01",X"00",X"C0",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"7F",X"3F",X"1E",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"00",X"00",
		X"FF",X"FF",X"FF",X"FB",X"F1",X"00",X"00",X"00",X"FF",X"FF",X"F7",X"E3",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"19",X"19",X"03",X"03",X"19",X"19",X"03",X"00",X"03",X"53",X"D8",X"03",X"D8",X"53",X"03",
		X"F8",X"48",X"EE",X"5F",X"89",X"FE",X"18",X"E8",X"FF",X"92",X"93",X"96",X"99",X"FF",X"33",X"D2",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",X"48",X"48",X"48",X"F8",X"58",X"58",X"58",X"48",
		X"92",X"92",X"92",X"BF",X"F2",X"F2",X"D2",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"68",X"F8",X"48",X"48",X"48",X"48",X"48",X"B2",X"92",X"9F",X"9A",X"BA",X"B2",X"92",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"58",X"58",X"58",X"48",X"68",X"68",X"F8",
		X"BF",X"F2",X"F2",X"D2",X"92",X"B2",X"92",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"48",X"48",X"48",X"FC",X"54",X"56",X"4A",X"9A",X"BA",X"B2",X"92",X"97",X"9E",X"9E",X"9A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"4A",X"FE",X"4A",X"4B",X"4D",X"4D",X"FF",X"48",
		X"92",X"97",X"9E",X"9E",X"9A",X"92",X"93",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"48",X"48",X"C8",X"C8",X"C8",X"48",X"48",X"97",X"96",X"92",X"92",X"93",X"93",X"FF",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"48",X"48",X"48",X"48",X"48",X"F8",X"48",X"F8",
		X"92",X"92",X"92",X"92",X"92",X"FF",X"92",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"78",X"98",X"F8",X"48",X"48",X"C8",X"C8",X"92",X"DE",X"96",X"F7",X"92",X"92",X"92",X"93",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"48",X"48",X"48",X"C8",X"C8",X"C8",X"48",
		X"93",X"FF",X"92",X"92",X"92",X"93",X"93",X"FF",X"00",X"03",X"02",X"02",X"02",X"02",X"02",X"03",
		X"48",X"FC",X"54",X"54",X"4C",X"48",X"F8",X"48",X"92",X"97",X"9E",X"9E",X"9A",X"92",X"BF",X"F2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"58",X"58",X"F8",X"48",X"48",X"48",X"48",
		X"F2",X"D2",X"92",X"9F",X"9A",X"BA",X"B2",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"F8",X"48",X"F8",X"48",X"C8",X"C8",X"C8",X"48",X"FF",X"92",X"FF",X"92",X"9F",X"90",X"9C",X"9D",
		X"02",X"02",X"04",X"04",X"04",X"04",X"04",X"04",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",
		X"92",X"92",X"92",X"AA",X"AA",X"AA",X"92",X"92",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",
		X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"48",X"48",X"48",X"F8",X"48",X"F8",X"F8",
		X"92",X"92",X"92",X"92",X"FF",X"92",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
